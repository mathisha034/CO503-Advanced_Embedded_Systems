// SoC.v

// Generated using ACDS version 13.1 162 at 2025.12.22.21:27:32

`timescale 1 ps / 1 ps
module SoC (
		input  wire        clk_clk,                            //                         clk.clk
		input  wire        reset_reset_n,                      //                       reset.reset_n
		output wire [12:0] sdram_addr,                         //                       sdram.addr
		output wire [1:0]  sdram_ba,                           //                            .ba
		output wire        sdram_cas_n,                        //                            .cas_n
		output wire        sdram_cke,                          //                            .cke
		output wire        sdram_cs_n,                         //                            .cs_n
		inout  wire [31:0] sdram_dq,                           //                            .dq
		output wire [3:0]  sdram_dqm,                          //                            .dqm
		output wire        sdram_ras_n,                        //                            .ras_n
		output wire        sdram_we_n,                         //                            .we_n
		output wire [7:0]  led_out_external_connection_export, // led_out_external_connection.export
		output wire        pll_c2_clk,                         //                      pll_c2.clk
		input  wire        pll_areset_conduit_export,          //          pll_areset_conduit.export
		output wire        pll_locked_conduit_export,          //          pll_locked_conduit.export
		output wire        pll_phasedone_conduit_export        //       pll_phasedone_conduit.export
	);

	wire         pll_c1_clk;                                                             // pll:c1 -> [irq_synchronizer:receiver_clk, mm_clock_crossing_bridge:m0_clk, mm_interconnect_1:pll_c1_clk, rst_controller_001:clk, sysid:clock, timer:clk]
	wire         pll_c0_clk;                                                             // pll:c0 -> [cpu:clk, irq_mapper:clk, irq_synchronizer:sender_clk, jtag_uart:clk, led_out:clk, mm_clock_crossing_bridge:s0_clk, mm_interconnect_0:pll_c0_clk, rst_controller:clk, sdram_controller:clk]
	wire  [31:0] cpu_custom_instruction_master_result;                                   // cpu_custom_instruction_master_translator:ci_slave_result -> cpu:E_ci_result
	wire   [4:0] cpu_custom_instruction_master_b;                                        // cpu:D_ci_b -> cpu_custom_instruction_master_translator:ci_slave_b
	wire   [4:0] cpu_custom_instruction_master_c;                                        // cpu:D_ci_c -> cpu_custom_instruction_master_translator:ci_slave_c
	wire         cpu_custom_instruction_master_done;                                     // cpu_custom_instruction_master_translator:ci_slave_multi_done -> cpu:E_ci_multi_done
	wire         cpu_custom_instruction_master_clk_en;                                   // cpu:E_ci_multi_clk_en -> cpu_custom_instruction_master_translator:ci_slave_multi_clken
	wire   [4:0] cpu_custom_instruction_master_a;                                        // cpu:D_ci_a -> cpu_custom_instruction_master_translator:ci_slave_a
	wire   [7:0] cpu_custom_instruction_master_n;                                        // cpu:D_ci_n -> cpu_custom_instruction_master_translator:ci_slave_n
	wire         cpu_custom_instruction_master_writerc;                                  // cpu:D_ci_writerc -> cpu_custom_instruction_master_translator:ci_slave_writerc
	wire         cpu_custom_instruction_master_clk;                                      // cpu:E_ci_multi_clock -> cpu_custom_instruction_master_translator:ci_slave_multi_clk
	wire         cpu_custom_instruction_master_reset_req;                                // cpu:E_ci_multi_reset_req -> cpu_custom_instruction_master_translator:ci_slave_multi_reset_req
	wire         cpu_custom_instruction_master_start;                                    // cpu:E_ci_multi_start -> cpu_custom_instruction_master_translator:ci_slave_multi_start
	wire  [31:0] cpu_custom_instruction_master_dataa;                                    // cpu:E_ci_dataa -> cpu_custom_instruction_master_translator:ci_slave_dataa
	wire         cpu_custom_instruction_master_readra;                                   // cpu:D_ci_readra -> cpu_custom_instruction_master_translator:ci_slave_readra
	wire         cpu_custom_instruction_master_reset;                                    // cpu:E_ci_multi_reset -> cpu_custom_instruction_master_translator:ci_slave_multi_reset
	wire  [31:0] cpu_custom_instruction_master_datab;                                    // cpu:E_ci_datab -> cpu_custom_instruction_master_translator:ci_slave_datab
	wire         cpu_custom_instruction_master_readrb;                                   // cpu:D_ci_readrb -> cpu_custom_instruction_master_translator:ci_slave_readrb
	wire  [31:0] cpu_custom_instruction_master_translator_multi_ci_master_result;        // cpu_custom_instruction_master_multi_xconnect:ci_slave_result -> cpu_custom_instruction_master_translator:multi_ci_master_result
	wire   [4:0] cpu_custom_instruction_master_translator_multi_ci_master_b;             // cpu_custom_instruction_master_translator:multi_ci_master_b -> cpu_custom_instruction_master_multi_xconnect:ci_slave_b
	wire   [4:0] cpu_custom_instruction_master_translator_multi_ci_master_c;             // cpu_custom_instruction_master_translator:multi_ci_master_c -> cpu_custom_instruction_master_multi_xconnect:ci_slave_c
	wire   [4:0] cpu_custom_instruction_master_translator_multi_ci_master_a;             // cpu_custom_instruction_master_translator:multi_ci_master_a -> cpu_custom_instruction_master_multi_xconnect:ci_slave_a
	wire         cpu_custom_instruction_master_translator_multi_ci_master_clk_en;        // cpu_custom_instruction_master_translator:multi_ci_master_clken -> cpu_custom_instruction_master_multi_xconnect:ci_slave_clken
	wire         cpu_custom_instruction_master_translator_multi_ci_master_done;          // cpu_custom_instruction_master_multi_xconnect:ci_slave_done -> cpu_custom_instruction_master_translator:multi_ci_master_done
	wire   [7:0] cpu_custom_instruction_master_translator_multi_ci_master_n;             // cpu_custom_instruction_master_translator:multi_ci_master_n -> cpu_custom_instruction_master_multi_xconnect:ci_slave_n
	wire         cpu_custom_instruction_master_translator_multi_ci_master_writerc;       // cpu_custom_instruction_master_translator:multi_ci_master_writerc -> cpu_custom_instruction_master_multi_xconnect:ci_slave_writerc
	wire         cpu_custom_instruction_master_translator_multi_ci_master_clk;           // cpu_custom_instruction_master_translator:multi_ci_master_clk -> cpu_custom_instruction_master_multi_xconnect:ci_slave_clk
	wire         cpu_custom_instruction_master_translator_multi_ci_master_reset_req;     // cpu_custom_instruction_master_translator:multi_ci_master_reset_req -> cpu_custom_instruction_master_multi_xconnect:ci_slave_reset_req
	wire         cpu_custom_instruction_master_translator_multi_ci_master_start;         // cpu_custom_instruction_master_translator:multi_ci_master_start -> cpu_custom_instruction_master_multi_xconnect:ci_slave_start
	wire  [31:0] cpu_custom_instruction_master_translator_multi_ci_master_dataa;         // cpu_custom_instruction_master_translator:multi_ci_master_dataa -> cpu_custom_instruction_master_multi_xconnect:ci_slave_dataa
	wire         cpu_custom_instruction_master_translator_multi_ci_master_readra;        // cpu_custom_instruction_master_translator:multi_ci_master_readra -> cpu_custom_instruction_master_multi_xconnect:ci_slave_readra
	wire         cpu_custom_instruction_master_translator_multi_ci_master_reset;         // cpu_custom_instruction_master_translator:multi_ci_master_reset -> cpu_custom_instruction_master_multi_xconnect:ci_slave_reset
	wire  [31:0] cpu_custom_instruction_master_translator_multi_ci_master_datab;         // cpu_custom_instruction_master_translator:multi_ci_master_datab -> cpu_custom_instruction_master_multi_xconnect:ci_slave_datab
	wire         cpu_custom_instruction_master_translator_multi_ci_master_readrb;        // cpu_custom_instruction_master_translator:multi_ci_master_readrb -> cpu_custom_instruction_master_multi_xconnect:ci_slave_readrb
	wire  [31:0] cpu_custom_instruction_master_multi_xconnect_ci_master0_result;         // cpu_custom_instruction_master_multi_slave_translator0:ci_slave_result -> cpu_custom_instruction_master_multi_xconnect:ci_master0_result
	wire   [4:0] cpu_custom_instruction_master_multi_xconnect_ci_master0_b;              // cpu_custom_instruction_master_multi_xconnect:ci_master0_b -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_b
	wire   [4:0] cpu_custom_instruction_master_multi_xconnect_ci_master0_c;              // cpu_custom_instruction_master_multi_xconnect:ci_master0_c -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_c
	wire         cpu_custom_instruction_master_multi_xconnect_ci_master0_done;           // cpu_custom_instruction_master_multi_slave_translator0:ci_slave_done -> cpu_custom_instruction_master_multi_xconnect:ci_master0_done
	wire         cpu_custom_instruction_master_multi_xconnect_ci_master0_clk_en;         // cpu_custom_instruction_master_multi_xconnect:ci_master0_clken -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_clken
	wire   [4:0] cpu_custom_instruction_master_multi_xconnect_ci_master0_a;              // cpu_custom_instruction_master_multi_xconnect:ci_master0_a -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_a
	wire   [7:0] cpu_custom_instruction_master_multi_xconnect_ci_master0_n;              // cpu_custom_instruction_master_multi_xconnect:ci_master0_n -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_n
	wire         cpu_custom_instruction_master_multi_xconnect_ci_master0_writerc;        // cpu_custom_instruction_master_multi_xconnect:ci_master0_writerc -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_writerc
	wire  [31:0] cpu_custom_instruction_master_multi_xconnect_ci_master0_ipending;       // cpu_custom_instruction_master_multi_xconnect:ci_master0_ipending -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_ipending
	wire         cpu_custom_instruction_master_multi_xconnect_ci_master0_clk;            // cpu_custom_instruction_master_multi_xconnect:ci_master0_clk -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_clk
	wire         cpu_custom_instruction_master_multi_xconnect_ci_master0_reset_req;      // cpu_custom_instruction_master_multi_xconnect:ci_master0_reset_req -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_reset_req
	wire         cpu_custom_instruction_master_multi_xconnect_ci_master0_start;          // cpu_custom_instruction_master_multi_xconnect:ci_master0_start -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_start
	wire  [31:0] cpu_custom_instruction_master_multi_xconnect_ci_master0_dataa;          // cpu_custom_instruction_master_multi_xconnect:ci_master0_dataa -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_dataa
	wire         cpu_custom_instruction_master_multi_xconnect_ci_master0_readra;         // cpu_custom_instruction_master_multi_xconnect:ci_master0_readra -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_readra
	wire         cpu_custom_instruction_master_multi_xconnect_ci_master0_reset;          // cpu_custom_instruction_master_multi_xconnect:ci_master0_reset -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_reset
	wire  [31:0] cpu_custom_instruction_master_multi_xconnect_ci_master0_datab;          // cpu_custom_instruction_master_multi_xconnect:ci_master0_datab -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_datab
	wire         cpu_custom_instruction_master_multi_xconnect_ci_master0_readrb;         // cpu_custom_instruction_master_multi_xconnect:ci_master0_readrb -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_readrb
	wire         cpu_custom_instruction_master_multi_xconnect_ci_master0_estatus;        // cpu_custom_instruction_master_multi_xconnect:ci_master0_estatus -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_estatus
	wire  [31:0] cpu_custom_instruction_master_multi_slave_translator0_ci_master_result; // CRC_0:result -> cpu_custom_instruction_master_multi_slave_translator0:ci_master_result
	wire         cpu_custom_instruction_master_multi_slave_translator0_ci_master_start;  // cpu_custom_instruction_master_multi_slave_translator0:ci_master_start -> CRC_0:start
	wire  [31:0] cpu_custom_instruction_master_multi_slave_translator0_ci_master_dataa;  // cpu_custom_instruction_master_multi_slave_translator0:ci_master_dataa -> CRC_0:dataa
	wire         cpu_custom_instruction_master_multi_slave_translator0_ci_master_done;   // CRC_0:done -> cpu_custom_instruction_master_multi_slave_translator0:ci_master_done
	wire         cpu_custom_instruction_master_multi_slave_translator0_ci_master_clk_en; // cpu_custom_instruction_master_multi_slave_translator0:ci_master_clken -> CRC_0:clk_en
	wire   [2:0] cpu_custom_instruction_master_multi_slave_translator0_ci_master_n;      // cpu_custom_instruction_master_multi_slave_translator0:ci_master_n -> CRC_0:n
	wire         cpu_custom_instruction_master_multi_slave_translator0_ci_master_reset;  // cpu_custom_instruction_master_multi_slave_translator0:ci_master_reset -> CRC_0:reset
	wire         cpu_custom_instruction_master_multi_slave_translator0_ci_master_clk;    // cpu_custom_instruction_master_multi_slave_translator0:ci_master_clk -> CRC_0:clk
	wire         mm_interconnect_0_cpu_jtag_debug_module_waitrequest;                    // cpu:jtag_debug_module_waitrequest -> mm_interconnect_0:cpu_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_cpu_jtag_debug_module_writedata;                      // mm_interconnect_0:cpu_jtag_debug_module_writedata -> cpu:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_cpu_jtag_debug_module_address;                        // mm_interconnect_0:cpu_jtag_debug_module_address -> cpu:jtag_debug_module_address
	wire         mm_interconnect_0_cpu_jtag_debug_module_write;                          // mm_interconnect_0:cpu_jtag_debug_module_write -> cpu:jtag_debug_module_write
	wire         mm_interconnect_0_cpu_jtag_debug_module_read;                           // mm_interconnect_0:cpu_jtag_debug_module_read -> cpu:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_cpu_jtag_debug_module_readdata;                       // cpu:jtag_debug_module_readdata -> mm_interconnect_0:cpu_jtag_debug_module_readdata
	wire         mm_interconnect_0_cpu_jtag_debug_module_debugaccess;                    // mm_interconnect_0:cpu_jtag_debug_module_debugaccess -> cpu:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_cpu_jtag_debug_module_byteenable;                     // mm_interconnect_0:cpu_jtag_debug_module_byteenable -> cpu:jtag_debug_module_byteenable
	wire  [31:0] mm_interconnect_0_pll_pll_slave_writedata;                              // mm_interconnect_0:pll_pll_slave_writedata -> pll:writedata
	wire   [1:0] mm_interconnect_0_pll_pll_slave_address;                                // mm_interconnect_0:pll_pll_slave_address -> pll:address
	wire         mm_interconnect_0_pll_pll_slave_write;                                  // mm_interconnect_0:pll_pll_slave_write -> pll:write
	wire         mm_interconnect_0_pll_pll_slave_read;                                   // mm_interconnect_0:pll_pll_slave_read -> pll:read
	wire  [31:0] mm_interconnect_0_pll_pll_slave_readdata;                               // pll:readdata -> mm_interconnect_0:pll_pll_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;              // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;                // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;                  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;               // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;                    // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;                     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;                 // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         cpu_data_master_waitrequest;                                            // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire  [31:0] cpu_data_master_writedata;                                              // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [27:0] cpu_data_master_address;                                                // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire         cpu_data_master_write;                                                  // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire         cpu_data_master_read;                                                   // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire  [31:0] cpu_data_master_readdata;                                               // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_debugaccess;                                            // cpu:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire   [3:0] cpu_data_master_byteenable;                                             // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire         cpu_instruction_master_waitrequest;                                     // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [27:0] cpu_instruction_master_address;                                         // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                                            // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire  [31:0] cpu_instruction_master_readdata;                                        // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire  [31:0] mm_interconnect_0_led_out_s1_writedata;                                 // mm_interconnect_0:led_out_s1_writedata -> led_out:writedata
	wire   [1:0] mm_interconnect_0_led_out_s1_address;                                   // mm_interconnect_0:led_out_s1_address -> led_out:address
	wire         mm_interconnect_0_led_out_s1_chipselect;                                // mm_interconnect_0:led_out_s1_chipselect -> led_out:chipselect
	wire         mm_interconnect_0_led_out_s1_write;                                     // mm_interconnect_0:led_out_s1_write -> led_out:write_n
	wire  [31:0] mm_interconnect_0_led_out_s1_readdata;                                  // led_out:readdata -> mm_interconnect_0:led_out_s1_readdata
	wire         mm_interconnect_0_sdram_controller_s1_waitrequest;                      // sdram_controller:za_waitrequest -> mm_interconnect_0:sdram_controller_s1_waitrequest
	wire  [31:0] mm_interconnect_0_sdram_controller_s1_writedata;                        // mm_interconnect_0:sdram_controller_s1_writedata -> sdram_controller:az_data
	wire  [24:0] mm_interconnect_0_sdram_controller_s1_address;                          // mm_interconnect_0:sdram_controller_s1_address -> sdram_controller:az_addr
	wire         mm_interconnect_0_sdram_controller_s1_chipselect;                       // mm_interconnect_0:sdram_controller_s1_chipselect -> sdram_controller:az_cs
	wire         mm_interconnect_0_sdram_controller_s1_write;                            // mm_interconnect_0:sdram_controller_s1_write -> sdram_controller:az_wr_n
	wire         mm_interconnect_0_sdram_controller_s1_read;                             // mm_interconnect_0:sdram_controller_s1_read -> sdram_controller:az_rd_n
	wire  [31:0] mm_interconnect_0_sdram_controller_s1_readdata;                         // sdram_controller:za_data -> mm_interconnect_0:sdram_controller_s1_readdata
	wire         mm_interconnect_0_sdram_controller_s1_readdatavalid;                    // sdram_controller:za_valid -> mm_interconnect_0:sdram_controller_s1_readdatavalid
	wire   [3:0] mm_interconnect_0_sdram_controller_s1_byteenable;                       // mm_interconnect_0:sdram_controller_s1_byteenable -> sdram_controller:az_be_n
	wire         mm_interconnect_0_mm_clock_crossing_bridge_s0_waitrequest;              // mm_clock_crossing_bridge:s0_waitrequest -> mm_interconnect_0:mm_clock_crossing_bridge_s0_waitrequest
	wire   [0:0] mm_interconnect_0_mm_clock_crossing_bridge_s0_burstcount;               // mm_interconnect_0:mm_clock_crossing_bridge_s0_burstcount -> mm_clock_crossing_bridge:s0_burstcount
	wire  [31:0] mm_interconnect_0_mm_clock_crossing_bridge_s0_writedata;                // mm_interconnect_0:mm_clock_crossing_bridge_s0_writedata -> mm_clock_crossing_bridge:s0_writedata
	wire   [9:0] mm_interconnect_0_mm_clock_crossing_bridge_s0_address;                  // mm_interconnect_0:mm_clock_crossing_bridge_s0_address -> mm_clock_crossing_bridge:s0_address
	wire         mm_interconnect_0_mm_clock_crossing_bridge_s0_write;                    // mm_interconnect_0:mm_clock_crossing_bridge_s0_write -> mm_clock_crossing_bridge:s0_write
	wire         mm_interconnect_0_mm_clock_crossing_bridge_s0_read;                     // mm_interconnect_0:mm_clock_crossing_bridge_s0_read -> mm_clock_crossing_bridge:s0_read
	wire  [31:0] mm_interconnect_0_mm_clock_crossing_bridge_s0_readdata;                 // mm_clock_crossing_bridge:s0_readdata -> mm_interconnect_0:mm_clock_crossing_bridge_s0_readdata
	wire         mm_interconnect_0_mm_clock_crossing_bridge_s0_debugaccess;              // mm_interconnect_0:mm_clock_crossing_bridge_s0_debugaccess -> mm_clock_crossing_bridge:s0_debugaccess
	wire         mm_interconnect_0_mm_clock_crossing_bridge_s0_readdatavalid;            // mm_clock_crossing_bridge:s0_readdatavalid -> mm_interconnect_0:mm_clock_crossing_bridge_s0_readdatavalid
	wire   [3:0] mm_interconnect_0_mm_clock_crossing_bridge_s0_byteenable;               // mm_interconnect_0:mm_clock_crossing_bridge_s0_byteenable -> mm_clock_crossing_bridge:s0_byteenable
	wire   [0:0] mm_interconnect_1_sysid_control_slave_address;                          // mm_interconnect_1:sysid_control_slave_address -> sysid:address
	wire  [31:0] mm_interconnect_1_sysid_control_slave_readdata;                         // sysid:readdata -> mm_interconnect_1:sysid_control_slave_readdata
	wire   [0:0] mm_clock_crossing_bridge_m0_burstcount;                                 // mm_clock_crossing_bridge:m0_burstcount -> mm_interconnect_1:mm_clock_crossing_bridge_m0_burstcount
	wire         mm_clock_crossing_bridge_m0_waitrequest;                                // mm_interconnect_1:mm_clock_crossing_bridge_m0_waitrequest -> mm_clock_crossing_bridge:m0_waitrequest
	wire   [9:0] mm_clock_crossing_bridge_m0_address;                                    // mm_clock_crossing_bridge:m0_address -> mm_interconnect_1:mm_clock_crossing_bridge_m0_address
	wire  [31:0] mm_clock_crossing_bridge_m0_writedata;                                  // mm_clock_crossing_bridge:m0_writedata -> mm_interconnect_1:mm_clock_crossing_bridge_m0_writedata
	wire         mm_clock_crossing_bridge_m0_write;                                      // mm_clock_crossing_bridge:m0_write -> mm_interconnect_1:mm_clock_crossing_bridge_m0_write
	wire         mm_clock_crossing_bridge_m0_read;                                       // mm_clock_crossing_bridge:m0_read -> mm_interconnect_1:mm_clock_crossing_bridge_m0_read
	wire  [31:0] mm_clock_crossing_bridge_m0_readdata;                                   // mm_interconnect_1:mm_clock_crossing_bridge_m0_readdata -> mm_clock_crossing_bridge:m0_readdata
	wire         mm_clock_crossing_bridge_m0_debugaccess;                                // mm_clock_crossing_bridge:m0_debugaccess -> mm_interconnect_1:mm_clock_crossing_bridge_m0_debugaccess
	wire   [3:0] mm_clock_crossing_bridge_m0_byteenable;                                 // mm_clock_crossing_bridge:m0_byteenable -> mm_interconnect_1:mm_clock_crossing_bridge_m0_byteenable
	wire         mm_clock_crossing_bridge_m0_readdatavalid;                              // mm_interconnect_1:mm_clock_crossing_bridge_m0_readdatavalid -> mm_clock_crossing_bridge:m0_readdatavalid
	wire  [15:0] mm_interconnect_1_timer_s1_writedata;                                   // mm_interconnect_1:timer_s1_writedata -> timer:writedata
	wire   [2:0] mm_interconnect_1_timer_s1_address;                                     // mm_interconnect_1:timer_s1_address -> timer:address
	wire         mm_interconnect_1_timer_s1_chipselect;                                  // mm_interconnect_1:timer_s1_chipselect -> timer:chipselect
	wire         mm_interconnect_1_timer_s1_write;                                       // mm_interconnect_1:timer_s1_write -> timer:write_n
	wire  [15:0] mm_interconnect_1_timer_s1_readdata;                                    // timer:readdata -> mm_interconnect_1:timer_s1_readdata
	wire         irq_mapper_receiver1_irq;                                               // jtag_uart:av_irq -> irq_mapper:receiver1_irq
	wire  [31:0] cpu_d_irq_irq;                                                          // irq_mapper:sender_irq -> cpu:d_irq
	wire         irq_mapper_receiver0_irq;                                               // irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	wire   [0:0] irq_synchronizer_receiver_irq;                                          // timer:irq -> irq_synchronizer:receiver_irq
	wire         rst_controller_reset_out_reset;                                         // rst_controller:reset_out -> [cpu:reset_n, irq_mapper:reset, irq_synchronizer:sender_reset, jtag_uart:rst_n, led_out:reset_n, mm_clock_crossing_bridge:s0_reset, mm_interconnect_0:cpu_reset_n_reset_bridge_in_reset_reset, rst_translator:in_reset, sdram_controller:reset_n]
	wire         rst_controller_reset_out_reset_req;                                     // rst_controller:reset_req -> [cpu:reset_req, rst_translator:reset_req_in]
	wire         cpu_jtag_debug_module_reset_reset;                                      // cpu:jtag_debug_module_resetrequest -> [rst_controller:reset_in1, rst_controller_001:reset_in1, rst_controller_002:reset_in1]
	wire         rst_controller_001_reset_out_reset;                                     // rst_controller_001:reset_out -> [irq_synchronizer:receiver_reset, mm_clock_crossing_bridge:m0_reset, mm_interconnect_1:mm_clock_crossing_bridge_m0_reset_reset_bridge_in_reset_reset, sysid:reset_n, timer:reset_n]
	wire         rst_controller_002_reset_out_reset;                                     // rst_controller_002:reset_out -> [mm_interconnect_0:pll_inclk_interface_reset_reset_bridge_in_reset_reset, pll:reset]

	SoC_sdram_controller sdram_controller (
		.clk            (pll_c0_clk),                                          //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),                     // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_controller_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_controller_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_controller_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_controller_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_controller_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_controller_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_controller_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_controller_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_controller_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_addr),                                          //  wire.export
		.zs_ba          (sdram_ba),                                            //      .export
		.zs_cas_n       (sdram_cas_n),                                         //      .export
		.zs_cke         (sdram_cke),                                           //      .export
		.zs_cs_n        (sdram_cs_n),                                          //      .export
		.zs_dq          (sdram_dq),                                            //      .export
		.zs_dqm         (sdram_dqm),                                           //      .export
		.zs_ras_n       (sdram_ras_n),                                         //      .export
		.zs_we_n        (sdram_we_n)                                           //      .export
	);

	SoC_cpu cpu (
		.clk                                   (pll_c0_clk),                                          //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                     //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                  //                          .reset_req
		.d_address                             (cpu_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpu_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpu_data_master_read),                                //                          .read
		.d_readdata                            (cpu_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpu_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpu_data_master_write),                               //                          .write
		.d_writedata                           (cpu_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpu_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpu_instruction_master_read),                         //                          .read
		.i_readdata                            (cpu_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpu_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (cpu_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_cpu_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_cpu_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_cpu_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_cpu_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_cpu_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_cpu_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_cpu_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_cpu_jtag_debug_module_writedata),   //                          .writedata
		.E_ci_multi_done                       (cpu_custom_instruction_master_done),                  // custom_instruction_master.done
		.E_ci_multi_clk_en                     (cpu_custom_instruction_master_clk_en),                //                          .clk_en
		.E_ci_multi_start                      (cpu_custom_instruction_master_start),                 //                          .start
		.E_ci_result                           (cpu_custom_instruction_master_result),                //                          .result
		.D_ci_a                                (cpu_custom_instruction_master_a),                     //                          .a
		.D_ci_b                                (cpu_custom_instruction_master_b),                     //                          .b
		.D_ci_c                                (cpu_custom_instruction_master_c),                     //                          .c
		.D_ci_n                                (cpu_custom_instruction_master_n),                     //                          .n
		.D_ci_readra                           (cpu_custom_instruction_master_readra),                //                          .readra
		.D_ci_readrb                           (cpu_custom_instruction_master_readrb),                //                          .readrb
		.D_ci_writerc                          (cpu_custom_instruction_master_writerc),               //                          .writerc
		.E_ci_dataa                            (cpu_custom_instruction_master_dataa),                 //                          .dataa
		.E_ci_datab                            (cpu_custom_instruction_master_datab),                 //                          .datab
		.E_ci_multi_clock                      (cpu_custom_instruction_master_clk),                   //                          .clk
		.E_ci_multi_reset                      (cpu_custom_instruction_master_reset),                 //                          .reset
		.E_ci_multi_reset_req                  (cpu_custom_instruction_master_reset_req)              //                          .reset_req
	);

	SoC_jtag_uart jtag_uart (
		.clk            (pll_c0_clk),                                                //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                   //               irq.irq
	);

	SoC_timer timer (
		.clk        (pll_c1_clk),                            //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),   // reset.reset_n
		.address    (mm_interconnect_1_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_1_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_1_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_1_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_1_timer_s1_write),     //      .write_n
		.irq        (irq_synchronizer_receiver_irq)          //   irq.irq
	);

	SoC_sysid sysid (
		.clock    (pll_c1_clk),                                     //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),            //         reset.reset_n
		.readdata (mm_interconnect_1_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_1_sysid_control_slave_address)   //              .address
	);

	SoC_led_out led_out (
		.clk        (pll_c0_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_led_out_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_out_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_out_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_out_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_out_s1_readdata),   //                    .readdata
		.out_port   (led_out_external_connection_export)       // external_connection.export
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.ADDRESS_WIDTH       (10),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (4),
		.RESPONSE_FIFO_DEPTH (4),
		.MASTER_SYNC_DEPTH   (2),
		.SLAVE_SYNC_DEPTH    (2)
	) mm_clock_crossing_bridge (
		.m0_clk           (pll_c1_clk),                                                  //   m0_clk.clk
		.m0_reset         (rst_controller_001_reset_out_reset),                          // m0_reset.reset
		.s0_clk           (pll_c0_clk),                                                  //   s0_clk.clk
		.s0_reset         (rst_controller_reset_out_reset),                              // s0_reset.reset
		.s0_waitrequest   (mm_interconnect_0_mm_clock_crossing_bridge_s0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (mm_interconnect_0_mm_clock_crossing_bridge_s0_readdata),      //         .readdata
		.s0_readdatavalid (mm_interconnect_0_mm_clock_crossing_bridge_s0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (mm_interconnect_0_mm_clock_crossing_bridge_s0_burstcount),    //         .burstcount
		.s0_writedata     (mm_interconnect_0_mm_clock_crossing_bridge_s0_writedata),     //         .writedata
		.s0_address       (mm_interconnect_0_mm_clock_crossing_bridge_s0_address),       //         .address
		.s0_write         (mm_interconnect_0_mm_clock_crossing_bridge_s0_write),         //         .write
		.s0_read          (mm_interconnect_0_mm_clock_crossing_bridge_s0_read),          //         .read
		.s0_byteenable    (mm_interconnect_0_mm_clock_crossing_bridge_s0_byteenable),    //         .byteenable
		.s0_debugaccess   (mm_interconnect_0_mm_clock_crossing_bridge_s0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (mm_clock_crossing_bridge_m0_waitrequest),                     //       m0.waitrequest
		.m0_readdata      (mm_clock_crossing_bridge_m0_readdata),                        //         .readdata
		.m0_readdatavalid (mm_clock_crossing_bridge_m0_readdatavalid),                   //         .readdatavalid
		.m0_burstcount    (mm_clock_crossing_bridge_m0_burstcount),                      //         .burstcount
		.m0_writedata     (mm_clock_crossing_bridge_m0_writedata),                       //         .writedata
		.m0_address       (mm_clock_crossing_bridge_m0_address),                         //         .address
		.m0_write         (mm_clock_crossing_bridge_m0_write),                           //         .write
		.m0_read          (mm_clock_crossing_bridge_m0_read),                            //         .read
		.m0_byteenable    (mm_clock_crossing_bridge_m0_byteenable),                      //         .byteenable
		.m0_debugaccess   (mm_clock_crossing_bridge_m0_debugaccess)                      //         .debugaccess
	);

	SoC_pll pll (
		.clk       (clk_clk),                                   //       inclk_interface.clk
		.reset     (rst_controller_002_reset_out_reset),        // inclk_interface_reset.reset
		.read      (mm_interconnect_0_pll_pll_slave_read),      //             pll_slave.read
		.write     (mm_interconnect_0_pll_pll_slave_write),     //                      .write
		.address   (mm_interconnect_0_pll_pll_slave_address),   //                      .address
		.readdata  (mm_interconnect_0_pll_pll_slave_readdata),  //                      .readdata
		.writedata (mm_interconnect_0_pll_pll_slave_writedata), //                      .writedata
		.c0        (pll_c0_clk),                                //                    c0.clk
		.c1        (pll_c1_clk),                                //                    c1.clk
		.c2        (pll_c2_clk),                                //                    c2.clk
		.areset    (pll_areset_conduit_export),                 //        areset_conduit.export
		.locked    (pll_locked_conduit_export),                 //        locked_conduit.export
		.phasedone (pll_phasedone_conduit_export)               //     phasedone_conduit.export
	);

	CRC_Custom_Instruction #(
		.crc_width         (32),
		.polynomial_inital (34'b0011111111111111111111111111111111),
		.polynomial        (34'b0000000100110000010001110110110111),
		.reflected_input   (1),
		.reflected_output  (1),
		.xor_output        (34'b0011111111111111111111111111111111)
	) crc_0 (
		.clk    (cpu_custom_instruction_master_multi_slave_translator0_ci_master_clk),    // nios_custom_instruction_slave.clk
		.reset  (cpu_custom_instruction_master_multi_slave_translator0_ci_master_reset),  //                              .reset
		.dataa  (cpu_custom_instruction_master_multi_slave_translator0_ci_master_dataa),  //                              .dataa
		.n      (cpu_custom_instruction_master_multi_slave_translator0_ci_master_n),      //                              .n
		.clk_en (cpu_custom_instruction_master_multi_slave_translator0_ci_master_clk_en), //                              .clk_en
		.start  (cpu_custom_instruction_master_multi_slave_translator0_ci_master_start),  //                              .start
		.done   (cpu_custom_instruction_master_multi_slave_translator0_ci_master_done),   //                              .done
		.result (cpu_custom_instruction_master_multi_slave_translator0_ci_master_result)  //                              .result
	);

	altera_customins_master_translator #(
		.SHARED_COMB_AND_MULTI (1)
	) cpu_custom_instruction_master_translator (
		.ci_slave_dataa            (cpu_custom_instruction_master_dataa),                                //        ci_slave.dataa
		.ci_slave_datab            (cpu_custom_instruction_master_datab),                                //                .datab
		.ci_slave_result           (cpu_custom_instruction_master_result),                               //                .result
		.ci_slave_n                (cpu_custom_instruction_master_n),                                    //                .n
		.ci_slave_readra           (cpu_custom_instruction_master_readra),                               //                .readra
		.ci_slave_readrb           (cpu_custom_instruction_master_readrb),                               //                .readrb
		.ci_slave_writerc          (cpu_custom_instruction_master_writerc),                              //                .writerc
		.ci_slave_a                (cpu_custom_instruction_master_a),                                    //                .a
		.ci_slave_b                (cpu_custom_instruction_master_b),                                    //                .b
		.ci_slave_c                (cpu_custom_instruction_master_c),                                    //                .c
		.ci_slave_ipending         (),                                                                   //                .ipending
		.ci_slave_estatus          (),                                                                   //                .estatus
		.ci_slave_multi_clk        (cpu_custom_instruction_master_clk),                                  //                .clk
		.ci_slave_multi_reset      (cpu_custom_instruction_master_reset),                                //                .reset
		.ci_slave_multi_clken      (cpu_custom_instruction_master_clk_en),                               //                .clk_en
		.ci_slave_multi_reset_req  (cpu_custom_instruction_master_reset_req),                            //                .reset_req
		.ci_slave_multi_start      (cpu_custom_instruction_master_start),                                //                .start
		.ci_slave_multi_done       (cpu_custom_instruction_master_done),                                 //                .done
		.comb_ci_master_dataa      (),                                                                   //  comb_ci_master.dataa
		.comb_ci_master_datab      (),                                                                   //                .datab
		.comb_ci_master_result     (),                                                                   //                .result
		.comb_ci_master_n          (),                                                                   //                .n
		.comb_ci_master_readra     (),                                                                   //                .readra
		.comb_ci_master_readrb     (),                                                                   //                .readrb
		.comb_ci_master_writerc    (),                                                                   //                .writerc
		.comb_ci_master_a          (),                                                                   //                .a
		.comb_ci_master_b          (),                                                                   //                .b
		.comb_ci_master_c          (),                                                                   //                .c
		.comb_ci_master_ipending   (),                                                                   //                .ipending
		.comb_ci_master_estatus    (),                                                                   //                .estatus
		.multi_ci_master_clk       (cpu_custom_instruction_master_translator_multi_ci_master_clk),       // multi_ci_master.clk
		.multi_ci_master_reset     (cpu_custom_instruction_master_translator_multi_ci_master_reset),     //                .reset
		.multi_ci_master_clken     (cpu_custom_instruction_master_translator_multi_ci_master_clk_en),    //                .clk_en
		.multi_ci_master_reset_req (cpu_custom_instruction_master_translator_multi_ci_master_reset_req), //                .reset_req
		.multi_ci_master_start     (cpu_custom_instruction_master_translator_multi_ci_master_start),     //                .start
		.multi_ci_master_done      (cpu_custom_instruction_master_translator_multi_ci_master_done),      //                .done
		.multi_ci_master_dataa     (cpu_custom_instruction_master_translator_multi_ci_master_dataa),     //                .dataa
		.multi_ci_master_datab     (cpu_custom_instruction_master_translator_multi_ci_master_datab),     //                .datab
		.multi_ci_master_result    (cpu_custom_instruction_master_translator_multi_ci_master_result),    //                .result
		.multi_ci_master_n         (cpu_custom_instruction_master_translator_multi_ci_master_n),         //                .n
		.multi_ci_master_readra    (cpu_custom_instruction_master_translator_multi_ci_master_readra),    //                .readra
		.multi_ci_master_readrb    (cpu_custom_instruction_master_translator_multi_ci_master_readrb),    //                .readrb
		.multi_ci_master_writerc   (cpu_custom_instruction_master_translator_multi_ci_master_writerc),   //                .writerc
		.multi_ci_master_a         (cpu_custom_instruction_master_translator_multi_ci_master_a),         //                .a
		.multi_ci_master_b         (cpu_custom_instruction_master_translator_multi_ci_master_b),         //                .b
		.multi_ci_master_c         (cpu_custom_instruction_master_translator_multi_ci_master_c),         //                .c
		.ci_slave_multi_dataa      (32'b00000000000000000000000000000000),                               //     (terminated)
		.ci_slave_multi_datab      (32'b00000000000000000000000000000000),                               //     (terminated)
		.ci_slave_multi_result     (),                                                                   //     (terminated)
		.ci_slave_multi_n          (8'b00000000),                                                        //     (terminated)
		.ci_slave_multi_readra     (1'b0),                                                               //     (terminated)
		.ci_slave_multi_readrb     (1'b0),                                                               //     (terminated)
		.ci_slave_multi_writerc    (1'b0),                                                               //     (terminated)
		.ci_slave_multi_a          (5'b00000),                                                           //     (terminated)
		.ci_slave_multi_b          (5'b00000),                                                           //     (terminated)
		.ci_slave_multi_c          (5'b00000)                                                            //     (terminated)
	);

	SoC_cpu_custom_instruction_master_multi_xconnect cpu_custom_instruction_master_multi_xconnect (
		.ci_slave_dataa       (cpu_custom_instruction_master_translator_multi_ci_master_dataa),     //   ci_slave.dataa
		.ci_slave_datab       (cpu_custom_instruction_master_translator_multi_ci_master_datab),     //           .datab
		.ci_slave_result      (cpu_custom_instruction_master_translator_multi_ci_master_result),    //           .result
		.ci_slave_n           (cpu_custom_instruction_master_translator_multi_ci_master_n),         //           .n
		.ci_slave_readra      (cpu_custom_instruction_master_translator_multi_ci_master_readra),    //           .readra
		.ci_slave_readrb      (cpu_custom_instruction_master_translator_multi_ci_master_readrb),    //           .readrb
		.ci_slave_writerc     (cpu_custom_instruction_master_translator_multi_ci_master_writerc),   //           .writerc
		.ci_slave_a           (cpu_custom_instruction_master_translator_multi_ci_master_a),         //           .a
		.ci_slave_b           (cpu_custom_instruction_master_translator_multi_ci_master_b),         //           .b
		.ci_slave_c           (cpu_custom_instruction_master_translator_multi_ci_master_c),         //           .c
		.ci_slave_ipending    (),                                                                   //           .ipending
		.ci_slave_estatus     (),                                                                   //           .estatus
		.ci_slave_clk         (cpu_custom_instruction_master_translator_multi_ci_master_clk),       //           .clk
		.ci_slave_reset       (cpu_custom_instruction_master_translator_multi_ci_master_reset),     //           .reset
		.ci_slave_clken       (cpu_custom_instruction_master_translator_multi_ci_master_clk_en),    //           .clk_en
		.ci_slave_reset_req   (cpu_custom_instruction_master_translator_multi_ci_master_reset_req), //           .reset_req
		.ci_slave_start       (cpu_custom_instruction_master_translator_multi_ci_master_start),     //           .start
		.ci_slave_done        (cpu_custom_instruction_master_translator_multi_ci_master_done),      //           .done
		.ci_master0_dataa     (cpu_custom_instruction_master_multi_xconnect_ci_master0_dataa),      // ci_master0.dataa
		.ci_master0_datab     (cpu_custom_instruction_master_multi_xconnect_ci_master0_datab),      //           .datab
		.ci_master0_result    (cpu_custom_instruction_master_multi_xconnect_ci_master0_result),     //           .result
		.ci_master0_n         (cpu_custom_instruction_master_multi_xconnect_ci_master0_n),          //           .n
		.ci_master0_readra    (cpu_custom_instruction_master_multi_xconnect_ci_master0_readra),     //           .readra
		.ci_master0_readrb    (cpu_custom_instruction_master_multi_xconnect_ci_master0_readrb),     //           .readrb
		.ci_master0_writerc   (cpu_custom_instruction_master_multi_xconnect_ci_master0_writerc),    //           .writerc
		.ci_master0_a         (cpu_custom_instruction_master_multi_xconnect_ci_master0_a),          //           .a
		.ci_master0_b         (cpu_custom_instruction_master_multi_xconnect_ci_master0_b),          //           .b
		.ci_master0_c         (cpu_custom_instruction_master_multi_xconnect_ci_master0_c),          //           .c
		.ci_master0_ipending  (cpu_custom_instruction_master_multi_xconnect_ci_master0_ipending),   //           .ipending
		.ci_master0_estatus   (cpu_custom_instruction_master_multi_xconnect_ci_master0_estatus),    //           .estatus
		.ci_master0_clk       (cpu_custom_instruction_master_multi_xconnect_ci_master0_clk),        //           .clk
		.ci_master0_reset     (cpu_custom_instruction_master_multi_xconnect_ci_master0_reset),      //           .reset
		.ci_master0_clken     (cpu_custom_instruction_master_multi_xconnect_ci_master0_clk_en),     //           .clk_en
		.ci_master0_reset_req (cpu_custom_instruction_master_multi_xconnect_ci_master0_reset_req),  //           .reset_req
		.ci_master0_start     (cpu_custom_instruction_master_multi_xconnect_ci_master0_start),      //           .start
		.ci_master0_done      (cpu_custom_instruction_master_multi_xconnect_ci_master0_done)        //           .done
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (3),
		.USE_DONE         (1),
		.NUM_FIXED_CYCLES (0)
	) cpu_custom_instruction_master_multi_slave_translator0 (
		.ci_slave_dataa      (cpu_custom_instruction_master_multi_xconnect_ci_master0_dataa),          //  ci_slave.dataa
		.ci_slave_datab      (cpu_custom_instruction_master_multi_xconnect_ci_master0_datab),          //          .datab
		.ci_slave_result     (cpu_custom_instruction_master_multi_xconnect_ci_master0_result),         //          .result
		.ci_slave_n          (cpu_custom_instruction_master_multi_xconnect_ci_master0_n),              //          .n
		.ci_slave_readra     (cpu_custom_instruction_master_multi_xconnect_ci_master0_readra),         //          .readra
		.ci_slave_readrb     (cpu_custom_instruction_master_multi_xconnect_ci_master0_readrb),         //          .readrb
		.ci_slave_writerc    (cpu_custom_instruction_master_multi_xconnect_ci_master0_writerc),        //          .writerc
		.ci_slave_a          (cpu_custom_instruction_master_multi_xconnect_ci_master0_a),              //          .a
		.ci_slave_b          (cpu_custom_instruction_master_multi_xconnect_ci_master0_b),              //          .b
		.ci_slave_c          (cpu_custom_instruction_master_multi_xconnect_ci_master0_c),              //          .c
		.ci_slave_ipending   (cpu_custom_instruction_master_multi_xconnect_ci_master0_ipending),       //          .ipending
		.ci_slave_estatus    (cpu_custom_instruction_master_multi_xconnect_ci_master0_estatus),        //          .estatus
		.ci_slave_clk        (cpu_custom_instruction_master_multi_xconnect_ci_master0_clk),            //          .clk
		.ci_slave_clken      (cpu_custom_instruction_master_multi_xconnect_ci_master0_clk_en),         //          .clk_en
		.ci_slave_reset_req  (cpu_custom_instruction_master_multi_xconnect_ci_master0_reset_req),      //          .reset_req
		.ci_slave_reset      (cpu_custom_instruction_master_multi_xconnect_ci_master0_reset),          //          .reset
		.ci_slave_start      (cpu_custom_instruction_master_multi_xconnect_ci_master0_start),          //          .start
		.ci_slave_done       (cpu_custom_instruction_master_multi_xconnect_ci_master0_done),           //          .done
		.ci_master_dataa     (cpu_custom_instruction_master_multi_slave_translator0_ci_master_dataa),  // ci_master.dataa
		.ci_master_result    (cpu_custom_instruction_master_multi_slave_translator0_ci_master_result), //          .result
		.ci_master_n         (cpu_custom_instruction_master_multi_slave_translator0_ci_master_n),      //          .n
		.ci_master_clk       (cpu_custom_instruction_master_multi_slave_translator0_ci_master_clk),    //          .clk
		.ci_master_clken     (cpu_custom_instruction_master_multi_slave_translator0_ci_master_clk_en), //          .clk_en
		.ci_master_reset     (cpu_custom_instruction_master_multi_slave_translator0_ci_master_reset),  //          .reset
		.ci_master_start     (cpu_custom_instruction_master_multi_slave_translator0_ci_master_start),  //          .start
		.ci_master_done      (cpu_custom_instruction_master_multi_slave_translator0_ci_master_done),   //          .done
		.ci_master_datab     (),                                                                       // (terminated)
		.ci_master_readra    (),                                                                       // (terminated)
		.ci_master_readrb    (),                                                                       // (terminated)
		.ci_master_writerc   (),                                                                       // (terminated)
		.ci_master_a         (),                                                                       // (terminated)
		.ci_master_b         (),                                                                       // (terminated)
		.ci_master_c         (),                                                                       // (terminated)
		.ci_master_ipending  (),                                                                       // (terminated)
		.ci_master_estatus   (),                                                                       // (terminated)
		.ci_master_reset_req ()                                                                        // (terminated)
	);

	SoC_mm_interconnect_0 mm_interconnect_0 (
		.clock_clk_clk                                         (clk_clk),                                                     //                                       clock_clk.clk
		.pll_c0_clk                                            (pll_c0_clk),                                                  //                                          pll_c0.clk
		.cpu_reset_n_reset_bridge_in_reset_reset               (rst_controller_reset_out_reset),                              //               cpu_reset_n_reset_bridge_in_reset.reset
		.pll_inclk_interface_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                          // pll_inclk_interface_reset_reset_bridge_in_reset.reset
		.cpu_data_master_address                               (cpu_data_master_address),                                     //                                 cpu_data_master.address
		.cpu_data_master_waitrequest                           (cpu_data_master_waitrequest),                                 //                                                .waitrequest
		.cpu_data_master_byteenable                            (cpu_data_master_byteenable),                                  //                                                .byteenable
		.cpu_data_master_read                                  (cpu_data_master_read),                                        //                                                .read
		.cpu_data_master_readdata                              (cpu_data_master_readdata),                                    //                                                .readdata
		.cpu_data_master_write                                 (cpu_data_master_write),                                       //                                                .write
		.cpu_data_master_writedata                             (cpu_data_master_writedata),                                   //                                                .writedata
		.cpu_data_master_debugaccess                           (cpu_data_master_debugaccess),                                 //                                                .debugaccess
		.cpu_instruction_master_address                        (cpu_instruction_master_address),                              //                          cpu_instruction_master.address
		.cpu_instruction_master_waitrequest                    (cpu_instruction_master_waitrequest),                          //                                                .waitrequest
		.cpu_instruction_master_read                           (cpu_instruction_master_read),                                 //                                                .read
		.cpu_instruction_master_readdata                       (cpu_instruction_master_readdata),                             //                                                .readdata
		.cpu_jtag_debug_module_address                         (mm_interconnect_0_cpu_jtag_debug_module_address),             //                           cpu_jtag_debug_module.address
		.cpu_jtag_debug_module_write                           (mm_interconnect_0_cpu_jtag_debug_module_write),               //                                                .write
		.cpu_jtag_debug_module_read                            (mm_interconnect_0_cpu_jtag_debug_module_read),                //                                                .read
		.cpu_jtag_debug_module_readdata                        (mm_interconnect_0_cpu_jtag_debug_module_readdata),            //                                                .readdata
		.cpu_jtag_debug_module_writedata                       (mm_interconnect_0_cpu_jtag_debug_module_writedata),           //                                                .writedata
		.cpu_jtag_debug_module_byteenable                      (mm_interconnect_0_cpu_jtag_debug_module_byteenable),          //                                                .byteenable
		.cpu_jtag_debug_module_waitrequest                     (mm_interconnect_0_cpu_jtag_debug_module_waitrequest),         //                                                .waitrequest
		.cpu_jtag_debug_module_debugaccess                     (mm_interconnect_0_cpu_jtag_debug_module_debugaccess),         //                                                .debugaccess
		.jtag_uart_avalon_jtag_slave_address                   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),       //                     jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),         //                                                .write
		.jtag_uart_avalon_jtag_slave_read                      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),          //                                                .read
		.jtag_uart_avalon_jtag_slave_readdata                  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),      //                                                .readdata
		.jtag_uart_avalon_jtag_slave_writedata                 (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),     //                                                .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest               (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),   //                                                .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),    //                                                .chipselect
		.led_out_s1_address                                    (mm_interconnect_0_led_out_s1_address),                        //                                      led_out_s1.address
		.led_out_s1_write                                      (mm_interconnect_0_led_out_s1_write),                          //                                                .write
		.led_out_s1_readdata                                   (mm_interconnect_0_led_out_s1_readdata),                       //                                                .readdata
		.led_out_s1_writedata                                  (mm_interconnect_0_led_out_s1_writedata),                      //                                                .writedata
		.led_out_s1_chipselect                                 (mm_interconnect_0_led_out_s1_chipselect),                     //                                                .chipselect
		.mm_clock_crossing_bridge_s0_address                   (mm_interconnect_0_mm_clock_crossing_bridge_s0_address),       //                     mm_clock_crossing_bridge_s0.address
		.mm_clock_crossing_bridge_s0_write                     (mm_interconnect_0_mm_clock_crossing_bridge_s0_write),         //                                                .write
		.mm_clock_crossing_bridge_s0_read                      (mm_interconnect_0_mm_clock_crossing_bridge_s0_read),          //                                                .read
		.mm_clock_crossing_bridge_s0_readdata                  (mm_interconnect_0_mm_clock_crossing_bridge_s0_readdata),      //                                                .readdata
		.mm_clock_crossing_bridge_s0_writedata                 (mm_interconnect_0_mm_clock_crossing_bridge_s0_writedata),     //                                                .writedata
		.mm_clock_crossing_bridge_s0_burstcount                (mm_interconnect_0_mm_clock_crossing_bridge_s0_burstcount),    //                                                .burstcount
		.mm_clock_crossing_bridge_s0_byteenable                (mm_interconnect_0_mm_clock_crossing_bridge_s0_byteenable),    //                                                .byteenable
		.mm_clock_crossing_bridge_s0_readdatavalid             (mm_interconnect_0_mm_clock_crossing_bridge_s0_readdatavalid), //                                                .readdatavalid
		.mm_clock_crossing_bridge_s0_waitrequest               (mm_interconnect_0_mm_clock_crossing_bridge_s0_waitrequest),   //                                                .waitrequest
		.mm_clock_crossing_bridge_s0_debugaccess               (mm_interconnect_0_mm_clock_crossing_bridge_s0_debugaccess),   //                                                .debugaccess
		.pll_pll_slave_address                                 (mm_interconnect_0_pll_pll_slave_address),                     //                                   pll_pll_slave.address
		.pll_pll_slave_write                                   (mm_interconnect_0_pll_pll_slave_write),                       //                                                .write
		.pll_pll_slave_read                                    (mm_interconnect_0_pll_pll_slave_read),                        //                                                .read
		.pll_pll_slave_readdata                                (mm_interconnect_0_pll_pll_slave_readdata),                    //                                                .readdata
		.pll_pll_slave_writedata                               (mm_interconnect_0_pll_pll_slave_writedata),                   //                                                .writedata
		.sdram_controller_s1_address                           (mm_interconnect_0_sdram_controller_s1_address),               //                             sdram_controller_s1.address
		.sdram_controller_s1_write                             (mm_interconnect_0_sdram_controller_s1_write),                 //                                                .write
		.sdram_controller_s1_read                              (mm_interconnect_0_sdram_controller_s1_read),                  //                                                .read
		.sdram_controller_s1_readdata                          (mm_interconnect_0_sdram_controller_s1_readdata),              //                                                .readdata
		.sdram_controller_s1_writedata                         (mm_interconnect_0_sdram_controller_s1_writedata),             //                                                .writedata
		.sdram_controller_s1_byteenable                        (mm_interconnect_0_sdram_controller_s1_byteenable),            //                                                .byteenable
		.sdram_controller_s1_readdatavalid                     (mm_interconnect_0_sdram_controller_s1_readdatavalid),         //                                                .readdatavalid
		.sdram_controller_s1_waitrequest                       (mm_interconnect_0_sdram_controller_s1_waitrequest),           //                                                .waitrequest
		.sdram_controller_s1_chipselect                        (mm_interconnect_0_sdram_controller_s1_chipselect)             //                                                .chipselect
	);

	SoC_mm_interconnect_1 mm_interconnect_1 (
		.pll_c1_clk                                                    (pll_c1_clk),                                     //                                                  pll_c1.clk
		.mm_clock_crossing_bridge_m0_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),             // mm_clock_crossing_bridge_m0_reset_reset_bridge_in_reset.reset
		.mm_clock_crossing_bridge_m0_address                           (mm_clock_crossing_bridge_m0_address),            //                             mm_clock_crossing_bridge_m0.address
		.mm_clock_crossing_bridge_m0_waitrequest                       (mm_clock_crossing_bridge_m0_waitrequest),        //                                                        .waitrequest
		.mm_clock_crossing_bridge_m0_burstcount                        (mm_clock_crossing_bridge_m0_burstcount),         //                                                        .burstcount
		.mm_clock_crossing_bridge_m0_byteenable                        (mm_clock_crossing_bridge_m0_byteenable),         //                                                        .byteenable
		.mm_clock_crossing_bridge_m0_read                              (mm_clock_crossing_bridge_m0_read),               //                                                        .read
		.mm_clock_crossing_bridge_m0_readdata                          (mm_clock_crossing_bridge_m0_readdata),           //                                                        .readdata
		.mm_clock_crossing_bridge_m0_readdatavalid                     (mm_clock_crossing_bridge_m0_readdatavalid),      //                                                        .readdatavalid
		.mm_clock_crossing_bridge_m0_write                             (mm_clock_crossing_bridge_m0_write),              //                                                        .write
		.mm_clock_crossing_bridge_m0_writedata                         (mm_clock_crossing_bridge_m0_writedata),          //                                                        .writedata
		.mm_clock_crossing_bridge_m0_debugaccess                       (mm_clock_crossing_bridge_m0_debugaccess),        //                                                        .debugaccess
		.sysid_control_slave_address                                   (mm_interconnect_1_sysid_control_slave_address),  //                                     sysid_control_slave.address
		.sysid_control_slave_readdata                                  (mm_interconnect_1_sysid_control_slave_readdata), //                                                        .readdata
		.timer_s1_address                                              (mm_interconnect_1_timer_s1_address),             //                                                timer_s1.address
		.timer_s1_write                                                (mm_interconnect_1_timer_s1_write),               //                                                        .write
		.timer_s1_readdata                                             (mm_interconnect_1_timer_s1_readdata),            //                                                        .readdata
		.timer_s1_writedata                                            (mm_interconnect_1_timer_s1_writedata),           //                                                        .writedata
		.timer_s1_chipselect                                           (mm_interconnect_1_timer_s1_chipselect)           //                                                        .chipselect
	);

	SoC_irq_mapper irq_mapper (
		.clk           (pll_c0_clk),                     //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (cpu_d_irq_irq)                   //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (pll_c1_clk),                         //       receiver_clk.clk
		.sender_clk     (pll_c0_clk),                         //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver0_irq)            //             sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_jtag_debug_module_reset_reset),  // reset_in1.reset
		.clk            (pll_c0_clk),                         //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_jtag_debug_module_reset_reset),  // reset_in1.reset
		.clk            (pll_c1_clk),                         //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_jtag_debug_module_reset_reset),  // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule

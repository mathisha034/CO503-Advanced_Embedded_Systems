// MPSoC.v

// Generated using ACDS version 13.1 162 at 2025.12.24.16:25:56

`timescale 1 ps / 1 ps
module MPSoC (
		input  wire  reset_reset_n, // reset.reset_n
		input  wire  clk_clk        //   clk.clk
	);

	wire         cpu_1_jtag_debug_module_reset_reset;                         // cpu_1:jtag_debug_module_resetrequest -> [jtag_uart_1:rst_n, mm_interconnect_0:jtag_uart_1_reset_reset_bridge_in_reset_reset, rst_controller_002:reset_in1, rst_controller_003:reset_in1]
	wire         cpu_1_data_master_waitrequest;                               // mm_interconnect_0:cpu_1_data_master_waitrequest -> cpu_1:d_waitrequest
	wire  [31:0] cpu_1_data_master_writedata;                                 // cpu_1:d_writedata -> mm_interconnect_0:cpu_1_data_master_writedata
	wire  [18:0] cpu_1_data_master_address;                                   // cpu_1:d_address -> mm_interconnect_0:cpu_1_data_master_address
	wire         cpu_1_data_master_write;                                     // cpu_1:d_write -> mm_interconnect_0:cpu_1_data_master_write
	wire         cpu_1_data_master_read;                                      // cpu_1:d_read -> mm_interconnect_0:cpu_1_data_master_read
	wire  [31:0] cpu_1_data_master_readdata;                                  // mm_interconnect_0:cpu_1_data_master_readdata -> cpu_1:d_readdata
	wire         cpu_1_data_master_debugaccess;                               // cpu_1:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:cpu_1_data_master_debugaccess
	wire   [3:0] cpu_1_data_master_byteenable;                                // cpu_1:d_byteenable -> mm_interconnect_0:cpu_1_data_master_byteenable
	wire         mm_interconnect_0_cpu_0_jtag_debug_module_waitrequest;       // cpu_0:jtag_debug_module_waitrequest -> mm_interconnect_0:cpu_0_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_cpu_0_jtag_debug_module_writedata;         // mm_interconnect_0:cpu_0_jtag_debug_module_writedata -> cpu_0:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_cpu_0_jtag_debug_module_address;           // mm_interconnect_0:cpu_0_jtag_debug_module_address -> cpu_0:jtag_debug_module_address
	wire         mm_interconnect_0_cpu_0_jtag_debug_module_write;             // mm_interconnect_0:cpu_0_jtag_debug_module_write -> cpu_0:jtag_debug_module_write
	wire         mm_interconnect_0_cpu_0_jtag_debug_module_read;              // mm_interconnect_0:cpu_0_jtag_debug_module_read -> cpu_0:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_cpu_0_jtag_debug_module_readdata;          // cpu_0:jtag_debug_module_readdata -> mm_interconnect_0:cpu_0_jtag_debug_module_readdata
	wire         mm_interconnect_0_cpu_0_jtag_debug_module_debugaccess;       // mm_interconnect_0:cpu_0_jtag_debug_module_debugaccess -> cpu_0:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_cpu_0_jtag_debug_module_byteenable;        // mm_interconnect_0:cpu_0_jtag_debug_module_byteenable -> cpu_0:jtag_debug_module_byteenable
	wire  [15:0] mm_interconnect_0_timer_1_s1_writedata;                      // mm_interconnect_0:timer_1_s1_writedata -> timer_1:writedata
	wire   [2:0] mm_interconnect_0_timer_1_s1_address;                        // mm_interconnect_0:timer_1_s1_address -> timer_1:address
	wire         mm_interconnect_0_timer_1_s1_chipselect;                     // mm_interconnect_0:timer_1_s1_chipselect -> timer_1:chipselect
	wire         mm_interconnect_0_timer_1_s1_write;                          // mm_interconnect_0:timer_1_s1_write -> timer_1:write_n
	wire  [15:0] mm_interconnect_0_timer_1_s1_readdata;                       // timer_1:readdata -> mm_interconnect_0:timer_1_s1_readdata
	wire   [0:0] mm_interconnect_0_sysid_0_control_slave_address;             // mm_interconnect_0:sysid_0_control_slave_address -> sysid_0:address
	wire  [31:0] mm_interconnect_0_sysid_0_control_slave_readdata;            // sysid_0:readdata -> mm_interconnect_0:sysid_0_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_1_control_slave_address;             // mm_interconnect_0:sysid_1_control_slave_address -> sysid_1:address
	wire  [31:0] mm_interconnect_0_sysid_1_control_slave_readdata;            // sysid_1:readdata -> mm_interconnect_0:sysid_1_control_slave_readdata
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                      // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                        // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_chipselect;                     // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire         mm_interconnect_0_timer_0_s1_write;                          // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                       // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire  [31:0] mm_interconnect_0_memory_shared_s1_writedata;                // mm_interconnect_0:memory_shared_s1_writedata -> memory_shared:writedata
	wire  [15:0] mm_interconnect_0_memory_shared_s1_address;                  // mm_interconnect_0:memory_shared_s1_address -> memory_shared:address
	wire         mm_interconnect_0_memory_shared_s1_chipselect;               // mm_interconnect_0:memory_shared_s1_chipselect -> memory_shared:chipselect
	wire         mm_interconnect_0_memory_shared_s1_clken;                    // mm_interconnect_0:memory_shared_s1_clken -> memory_shared:clken
	wire         mm_interconnect_0_memory_shared_s1_write;                    // mm_interconnect_0:memory_shared_s1_write -> memory_shared:write
	wire  [31:0] mm_interconnect_0_memory_shared_s1_readdata;                 // memory_shared:readdata -> mm_interconnect_0:memory_shared_s1_readdata
	wire   [3:0] mm_interconnect_0_memory_shared_s1_byteenable;               // mm_interconnect_0:memory_shared_s1_byteenable -> memory_shared:byteenable
	wire         mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_waitrequest; // jtag_uart_1:av_waitrequest -> mm_interconnect_0:jtag_uart_1_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_1_avalon_jtag_slave_writedata -> jtag_uart_1:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_1_avalon_jtag_slave_address -> jtag_uart_1:av_address
	wire         mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_1_avalon_jtag_slave_chipselect -> jtag_uart_1:av_chipselect
	wire         mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_1_avalon_jtag_slave_write -> jtag_uart_1:av_write_n
	wire         mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_1_avalon_jtag_slave_read -> jtag_uart_1:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_readdata;    // jtag_uart_1:av_readdata -> mm_interconnect_0:jtag_uart_1_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_cpu_1_jtag_debug_module_waitrequest;       // cpu_1:jtag_debug_module_waitrequest -> mm_interconnect_0:cpu_1_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_cpu_1_jtag_debug_module_writedata;         // mm_interconnect_0:cpu_1_jtag_debug_module_writedata -> cpu_1:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_cpu_1_jtag_debug_module_address;           // mm_interconnect_0:cpu_1_jtag_debug_module_address -> cpu_1:jtag_debug_module_address
	wire         mm_interconnect_0_cpu_1_jtag_debug_module_write;             // mm_interconnect_0:cpu_1_jtag_debug_module_write -> cpu_1:jtag_debug_module_write
	wire         mm_interconnect_0_cpu_1_jtag_debug_module_read;              // mm_interconnect_0:cpu_1_jtag_debug_module_read -> cpu_1:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_cpu_1_jtag_debug_module_readdata;          // cpu_1:jtag_debug_module_readdata -> mm_interconnect_0:cpu_1_jtag_debug_module_readdata
	wire         mm_interconnect_0_cpu_1_jtag_debug_module_debugaccess;       // mm_interconnect_0:cpu_1_jtag_debug_module_debugaccess -> cpu_1:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_cpu_1_jtag_debug_module_byteenable;        // mm_interconnect_0:cpu_1_jtag_debug_module_byteenable -> cpu_1:jtag_debug_module_byteenable
	wire         cpu_0_instruction_master_waitrequest;                        // mm_interconnect_0:cpu_0_instruction_master_waitrequest -> cpu_0:i_waitrequest
	wire  [18:0] cpu_0_instruction_master_address;                            // cpu_0:i_address -> mm_interconnect_0:cpu_0_instruction_master_address
	wire         cpu_0_instruction_master_read;                               // cpu_0:i_read -> mm_interconnect_0:cpu_0_instruction_master_read
	wire  [31:0] cpu_0_instruction_master_readdata;                           // mm_interconnect_0:cpu_0_instruction_master_readdata -> cpu_0:i_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         cpu_0_data_master_waitrequest;                               // mm_interconnect_0:cpu_0_data_master_waitrequest -> cpu_0:d_waitrequest
	wire  [31:0] cpu_0_data_master_writedata;                                 // cpu_0:d_writedata -> mm_interconnect_0:cpu_0_data_master_writedata
	wire  [18:0] cpu_0_data_master_address;                                   // cpu_0:d_address -> mm_interconnect_0:cpu_0_data_master_address
	wire         cpu_0_data_master_write;                                     // cpu_0:d_write -> mm_interconnect_0:cpu_0_data_master_write
	wire         cpu_0_data_master_read;                                      // cpu_0:d_read -> mm_interconnect_0:cpu_0_data_master_read
	wire  [31:0] cpu_0_data_master_readdata;                                  // mm_interconnect_0:cpu_0_data_master_readdata -> cpu_0:d_readdata
	wire         cpu_0_data_master_debugaccess;                               // cpu_0:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:cpu_0_data_master_debugaccess
	wire   [3:0] cpu_0_data_master_byteenable;                                // cpu_0:d_byteenable -> mm_interconnect_0:cpu_0_data_master_byteenable
	wire         cpu_1_instruction_master_waitrequest;                        // mm_interconnect_0:cpu_1_instruction_master_waitrequest -> cpu_1:i_waitrequest
	wire  [18:0] cpu_1_instruction_master_address;                            // cpu_1:i_address -> mm_interconnect_0:cpu_1_instruction_master_address
	wire         cpu_1_instruction_master_read;                               // cpu_1:i_read -> mm_interconnect_0:cpu_1_instruction_master_read
	wire  [31:0] cpu_1_instruction_master_readdata;                           // mm_interconnect_0:cpu_1_instruction_master_readdata -> cpu_1:i_readdata
	wire  [31:0] mm_interconnect_0_memory_0_s1_writedata;                     // mm_interconnect_0:memory_0_s1_writedata -> memory_0:writedata
	wire  [14:0] mm_interconnect_0_memory_0_s1_address;                       // mm_interconnect_0:memory_0_s1_address -> memory_0:address
	wire         mm_interconnect_0_memory_0_s1_chipselect;                    // mm_interconnect_0:memory_0_s1_chipselect -> memory_0:chipselect
	wire         mm_interconnect_0_memory_0_s1_clken;                         // mm_interconnect_0:memory_0_s1_clken -> memory_0:clken
	wire         mm_interconnect_0_memory_0_s1_write;                         // mm_interconnect_0:memory_0_s1_write -> memory_0:write
	wire  [31:0] mm_interconnect_0_memory_0_s1_readdata;                      // memory_0:readdata -> mm_interconnect_0:memory_0_s1_readdata
	wire   [3:0] mm_interconnect_0_memory_0_s1_byteenable;                    // mm_interconnect_0:memory_0_s1_byteenable -> memory_0:byteenable
	wire  [31:0] mm_interconnect_0_memory_1_s1_writedata;                     // mm_interconnect_0:memory_1_s1_writedata -> memory_1:writedata
	wire  [14:0] mm_interconnect_0_memory_1_s1_address;                       // mm_interconnect_0:memory_1_s1_address -> memory_1:address
	wire         mm_interconnect_0_memory_1_s1_chipselect;                    // mm_interconnect_0:memory_1_s1_chipselect -> memory_1:chipselect
	wire         mm_interconnect_0_memory_1_s1_clken;                         // mm_interconnect_0:memory_1_s1_clken -> memory_1:clken
	wire         mm_interconnect_0_memory_1_s1_write;                         // mm_interconnect_0:memory_1_s1_write -> memory_1:write
	wire  [31:0] mm_interconnect_0_memory_1_s1_readdata;                      // memory_1:readdata -> mm_interconnect_0:memory_1_s1_readdata
	wire   [3:0] mm_interconnect_0_memory_1_s1_byteenable;                    // mm_interconnect_0:memory_1_s1_byteenable -> memory_1:byteenable
	wire         irq_mapper_receiver0_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                    // timer_0:irq -> irq_mapper:receiver1_irq
	wire  [31:0] cpu_0_d_irq_irq;                                             // irq_mapper:sender_irq -> cpu_0:d_irq
	wire         irq_mapper_001_receiver0_irq;                                // timer_1:irq -> irq_mapper_001:receiver0_irq
	wire         irq_mapper_001_receiver1_irq;                                // jtag_uart_1:av_irq -> irq_mapper_001:receiver1_irq
	wire  [31:0] cpu_1_d_irq_irq;                                             // irq_mapper_001:sender_irq -> cpu_1:d_irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [jtag_uart_0:rst_n, memory_0:reset, mm_interconnect_0:memory_0_reset1_reset_bridge_in_reset_reset, rst_translator:in_reset, sysid_0:reset_n, timer_0:reset_n]
	wire         rst_controller_reset_out_reset_req;                          // rst_controller:reset_req -> [memory_0:reset_req, rst_translator:reset_req_in]
	wire         cpu_0_jtag_debug_module_reset_reset;                         // cpu_0:jtag_debug_module_resetrequest -> [rst_controller:reset_in1, rst_controller_003:reset_in2]
	wire         rst_controller_001_reset_out_reset;                          // rst_controller_001:reset_out -> [cpu_0:reset_n, cpu_1:reset_n, irq_mapper:reset, irq_mapper_001:reset, mm_interconnect_0:cpu_0_reset_n_reset_bridge_in_reset_reset, rst_translator_001:in_reset]
	wire         rst_controller_001_reset_out_reset_req;                      // rst_controller_001:reset_req -> [cpu_0:reset_req, cpu_1:reset_req, rst_translator_001:reset_req_in]
	wire         rst_controller_002_reset_out_reset;                          // rst_controller_002:reset_out -> [memory_1:reset, mm_interconnect_0:timer_1_reset_reset_bridge_in_reset_reset, rst_translator_002:in_reset, sysid_1:reset_n, timer_1:reset_n]
	wire         rst_controller_002_reset_out_reset_req;                      // rst_controller_002:reset_req -> [memory_1:reset_req, rst_translator_002:reset_req_in]
	wire         rst_controller_003_reset_out_reset;                          // rst_controller_003:reset_out -> [memory_shared:reset, mm_interconnect_0:memory_shared_reset1_reset_bridge_in_reset_reset]
	wire         rst_controller_003_reset_out_reset_req;                      // rst_controller_003:reset_req -> memory_shared:reset_req

	MPSoC_memory_0 memory_0 (
		.clk        (clk_clk),                                  //   clk1.clk
		.address    (mm_interconnect_0_memory_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_memory_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_memory_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_memory_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_memory_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_memory_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_memory_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),           // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)        //       .reset_req
	);

	MPSoC_cpu_0 cpu_0 (
		.clk                                   (clk_clk),                                               //                       clk.clk
		.reset_n                               (~rst_controller_001_reset_out_reset),                   //                   reset_n.reset_n
		.reset_req                             (rst_controller_001_reset_out_reset_req),                //                          .reset_req
		.d_address                             (cpu_0_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpu_0_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpu_0_data_master_read),                                //                          .read
		.d_readdata                            (cpu_0_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpu_0_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpu_0_data_master_write),                               //                          .write
		.d_writedata                           (cpu_0_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_0_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpu_0_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpu_0_instruction_master_read),                         //                          .read
		.i_readdata                            (cpu_0_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpu_0_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (cpu_0_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_0_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_cpu_0_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_cpu_0_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_cpu_0_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_cpu_0_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_cpu_0_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_cpu_0_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_cpu_0_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_cpu_0_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                       // custom_instruction_master.readra
	);

	MPSoC_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	MPSoC_timer_0 timer_0 (
		.clk        (clk_clk),                                 //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                 //   irq.irq
	);

	MPSoC_sysid_0 sysid_0 (
		.clock    (clk_clk),                                          //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                  //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_0_control_slave_address)   //              .address
	);

	MPSoC_memory_1 memory_1 (
		.clk        (clk_clk),                                  //   clk1.clk
		.address    (mm_interconnect_0_memory_1_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_memory_1_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_memory_1_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_memory_1_s1_write),      //       .write
		.readdata   (mm_interconnect_0_memory_1_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_memory_1_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_memory_1_s1_byteenable), //       .byteenable
		.reset      (rst_controller_002_reset_out_reset),       // reset1.reset
		.reset_req  (rst_controller_002_reset_out_reset_req)    //       .reset_req
	);

	MPSoC_cpu_1 cpu_1 (
		.clk                                   (clk_clk),                                               //                       clk.clk
		.reset_n                               (~rst_controller_001_reset_out_reset),                   //                   reset_n.reset_n
		.reset_req                             (rst_controller_001_reset_out_reset_req),                //                          .reset_req
		.d_address                             (cpu_1_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpu_1_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpu_1_data_master_read),                                //                          .read
		.d_readdata                            (cpu_1_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpu_1_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpu_1_data_master_write),                               //                          .write
		.d_writedata                           (cpu_1_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_1_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpu_1_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpu_1_instruction_master_read),                         //                          .read
		.i_readdata                            (cpu_1_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpu_1_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (cpu_1_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_1_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_cpu_1_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_cpu_1_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_cpu_1_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_cpu_1_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_cpu_1_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_cpu_1_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_cpu_1_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_cpu_1_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                       // custom_instruction_master.readra
	);

	MPSoC_jtag_uart_0 jtag_uart_1 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~cpu_1_jtag_debug_module_reset_reset),                        //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_001_receiver1_irq)                                 //               irq.irq
	);

	MPSoC_timer_0 timer_1 (
		.clk        (clk_clk),                                 //   clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),     // reset.reset_n
		.address    (mm_interconnect_0_timer_1_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_1_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_1_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_1_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_1_s1_write),     //      .write_n
		.irq        (irq_mapper_001_receiver0_irq)             //   irq.irq
	);

	MPSoC_sysid_0 sysid_1 (
		.clock    (clk_clk),                                          //           clk.clk
		.reset_n  (~rst_controller_002_reset_out_reset),              //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_1_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_1_control_slave_address)   //              .address
	);

	MPSoC_memory_shared memory_shared (
		.clk        (clk_clk),                                       //   clk1.clk
		.address    (mm_interconnect_0_memory_shared_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_memory_shared_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_memory_shared_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_memory_shared_s1_write),      //       .write
		.readdata   (mm_interconnect_0_memory_shared_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_memory_shared_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_memory_shared_s1_byteenable), //       .byteenable
		.reset      (rst_controller_003_reset_out_reset),            // reset1.reset
		.reset_req  (rst_controller_003_reset_out_reset_req)         //       .reset_req
	);

	MPSoC_mm_interconnect_0 mm_interconnect_0 (
		.clock_clk_clk                                    (clk_clk),                                                     //                                  clock_clk.clk
		.cpu_0_reset_n_reset_bridge_in_reset_reset        (rst_controller_001_reset_out_reset),                          //        cpu_0_reset_n_reset_bridge_in_reset.reset
		.jtag_uart_1_reset_reset_bridge_in_reset_reset    (cpu_1_jtag_debug_module_reset_reset),                         //    jtag_uart_1_reset_reset_bridge_in_reset.reset
		.memory_0_reset1_reset_bridge_in_reset_reset      (rst_controller_reset_out_reset),                              //      memory_0_reset1_reset_bridge_in_reset.reset
		.memory_shared_reset1_reset_bridge_in_reset_reset (rst_controller_003_reset_out_reset),                          // memory_shared_reset1_reset_bridge_in_reset.reset
		.timer_1_reset_reset_bridge_in_reset_reset        (rst_controller_002_reset_out_reset),                          //        timer_1_reset_reset_bridge_in_reset.reset
		.cpu_0_data_master_address                        (cpu_0_data_master_address),                                   //                          cpu_0_data_master.address
		.cpu_0_data_master_waitrequest                    (cpu_0_data_master_waitrequest),                               //                                           .waitrequest
		.cpu_0_data_master_byteenable                     (cpu_0_data_master_byteenable),                                //                                           .byteenable
		.cpu_0_data_master_read                           (cpu_0_data_master_read),                                      //                                           .read
		.cpu_0_data_master_readdata                       (cpu_0_data_master_readdata),                                  //                                           .readdata
		.cpu_0_data_master_write                          (cpu_0_data_master_write),                                     //                                           .write
		.cpu_0_data_master_writedata                      (cpu_0_data_master_writedata),                                 //                                           .writedata
		.cpu_0_data_master_debugaccess                    (cpu_0_data_master_debugaccess),                               //                                           .debugaccess
		.cpu_0_instruction_master_address                 (cpu_0_instruction_master_address),                            //                   cpu_0_instruction_master.address
		.cpu_0_instruction_master_waitrequest             (cpu_0_instruction_master_waitrequest),                        //                                           .waitrequest
		.cpu_0_instruction_master_read                    (cpu_0_instruction_master_read),                               //                                           .read
		.cpu_0_instruction_master_readdata                (cpu_0_instruction_master_readdata),                           //                                           .readdata
		.cpu_1_data_master_address                        (cpu_1_data_master_address),                                   //                          cpu_1_data_master.address
		.cpu_1_data_master_waitrequest                    (cpu_1_data_master_waitrequest),                               //                                           .waitrequest
		.cpu_1_data_master_byteenable                     (cpu_1_data_master_byteenable),                                //                                           .byteenable
		.cpu_1_data_master_read                           (cpu_1_data_master_read),                                      //                                           .read
		.cpu_1_data_master_readdata                       (cpu_1_data_master_readdata),                                  //                                           .readdata
		.cpu_1_data_master_write                          (cpu_1_data_master_write),                                     //                                           .write
		.cpu_1_data_master_writedata                      (cpu_1_data_master_writedata),                                 //                                           .writedata
		.cpu_1_data_master_debugaccess                    (cpu_1_data_master_debugaccess),                               //                                           .debugaccess
		.cpu_1_instruction_master_address                 (cpu_1_instruction_master_address),                            //                   cpu_1_instruction_master.address
		.cpu_1_instruction_master_waitrequest             (cpu_1_instruction_master_waitrequest),                        //                                           .waitrequest
		.cpu_1_instruction_master_read                    (cpu_1_instruction_master_read),                               //                                           .read
		.cpu_1_instruction_master_readdata                (cpu_1_instruction_master_readdata),                           //                                           .readdata
		.cpu_0_jtag_debug_module_address                  (mm_interconnect_0_cpu_0_jtag_debug_module_address),           //                    cpu_0_jtag_debug_module.address
		.cpu_0_jtag_debug_module_write                    (mm_interconnect_0_cpu_0_jtag_debug_module_write),             //                                           .write
		.cpu_0_jtag_debug_module_read                     (mm_interconnect_0_cpu_0_jtag_debug_module_read),              //                                           .read
		.cpu_0_jtag_debug_module_readdata                 (mm_interconnect_0_cpu_0_jtag_debug_module_readdata),          //                                           .readdata
		.cpu_0_jtag_debug_module_writedata                (mm_interconnect_0_cpu_0_jtag_debug_module_writedata),         //                                           .writedata
		.cpu_0_jtag_debug_module_byteenable               (mm_interconnect_0_cpu_0_jtag_debug_module_byteenable),        //                                           .byteenable
		.cpu_0_jtag_debug_module_waitrequest              (mm_interconnect_0_cpu_0_jtag_debug_module_waitrequest),       //                                           .waitrequest
		.cpu_0_jtag_debug_module_debugaccess              (mm_interconnect_0_cpu_0_jtag_debug_module_debugaccess),       //                                           .debugaccess
		.cpu_1_jtag_debug_module_address                  (mm_interconnect_0_cpu_1_jtag_debug_module_address),           //                    cpu_1_jtag_debug_module.address
		.cpu_1_jtag_debug_module_write                    (mm_interconnect_0_cpu_1_jtag_debug_module_write),             //                                           .write
		.cpu_1_jtag_debug_module_read                     (mm_interconnect_0_cpu_1_jtag_debug_module_read),              //                                           .read
		.cpu_1_jtag_debug_module_readdata                 (mm_interconnect_0_cpu_1_jtag_debug_module_readdata),          //                                           .readdata
		.cpu_1_jtag_debug_module_writedata                (mm_interconnect_0_cpu_1_jtag_debug_module_writedata),         //                                           .writedata
		.cpu_1_jtag_debug_module_byteenable               (mm_interconnect_0_cpu_1_jtag_debug_module_byteenable),        //                                           .byteenable
		.cpu_1_jtag_debug_module_waitrequest              (mm_interconnect_0_cpu_1_jtag_debug_module_waitrequest),       //                                           .waitrequest
		.cpu_1_jtag_debug_module_debugaccess              (mm_interconnect_0_cpu_1_jtag_debug_module_debugaccess),       //                                           .debugaccess
		.jtag_uart_0_avalon_jtag_slave_address            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //              jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write              (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                           .write
		.jtag_uart_0_avalon_jtag_slave_read               (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                           .read
		.jtag_uart_0_avalon_jtag_slave_readdata           (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                           .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                           .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                           .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                           .chipselect
		.jtag_uart_1_avalon_jtag_slave_address            (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_address),     //              jtag_uart_1_avalon_jtag_slave.address
		.jtag_uart_1_avalon_jtag_slave_write              (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_write),       //                                           .write
		.jtag_uart_1_avalon_jtag_slave_read               (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_read),        //                                           .read
		.jtag_uart_1_avalon_jtag_slave_readdata           (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_readdata),    //                                           .readdata
		.jtag_uart_1_avalon_jtag_slave_writedata          (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_writedata),   //                                           .writedata
		.jtag_uart_1_avalon_jtag_slave_waitrequest        (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_waitrequest), //                                           .waitrequest
		.jtag_uart_1_avalon_jtag_slave_chipselect         (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_chipselect),  //                                           .chipselect
		.memory_0_s1_address                              (mm_interconnect_0_memory_0_s1_address),                       //                                memory_0_s1.address
		.memory_0_s1_write                                (mm_interconnect_0_memory_0_s1_write),                         //                                           .write
		.memory_0_s1_readdata                             (mm_interconnect_0_memory_0_s1_readdata),                      //                                           .readdata
		.memory_0_s1_writedata                            (mm_interconnect_0_memory_0_s1_writedata),                     //                                           .writedata
		.memory_0_s1_byteenable                           (mm_interconnect_0_memory_0_s1_byteenable),                    //                                           .byteenable
		.memory_0_s1_chipselect                           (mm_interconnect_0_memory_0_s1_chipselect),                    //                                           .chipselect
		.memory_0_s1_clken                                (mm_interconnect_0_memory_0_s1_clken),                         //                                           .clken
		.memory_1_s1_address                              (mm_interconnect_0_memory_1_s1_address),                       //                                memory_1_s1.address
		.memory_1_s1_write                                (mm_interconnect_0_memory_1_s1_write),                         //                                           .write
		.memory_1_s1_readdata                             (mm_interconnect_0_memory_1_s1_readdata),                      //                                           .readdata
		.memory_1_s1_writedata                            (mm_interconnect_0_memory_1_s1_writedata),                     //                                           .writedata
		.memory_1_s1_byteenable                           (mm_interconnect_0_memory_1_s1_byteenable),                    //                                           .byteenable
		.memory_1_s1_chipselect                           (mm_interconnect_0_memory_1_s1_chipselect),                    //                                           .chipselect
		.memory_1_s1_clken                                (mm_interconnect_0_memory_1_s1_clken),                         //                                           .clken
		.memory_shared_s1_address                         (mm_interconnect_0_memory_shared_s1_address),                  //                           memory_shared_s1.address
		.memory_shared_s1_write                           (mm_interconnect_0_memory_shared_s1_write),                    //                                           .write
		.memory_shared_s1_readdata                        (mm_interconnect_0_memory_shared_s1_readdata),                 //                                           .readdata
		.memory_shared_s1_writedata                       (mm_interconnect_0_memory_shared_s1_writedata),                //                                           .writedata
		.memory_shared_s1_byteenable                      (mm_interconnect_0_memory_shared_s1_byteenable),               //                                           .byteenable
		.memory_shared_s1_chipselect                      (mm_interconnect_0_memory_shared_s1_chipselect),               //                                           .chipselect
		.memory_shared_s1_clken                           (mm_interconnect_0_memory_shared_s1_clken),                    //                                           .clken
		.sysid_0_control_slave_address                    (mm_interconnect_0_sysid_0_control_slave_address),             //                      sysid_0_control_slave.address
		.sysid_0_control_slave_readdata                   (mm_interconnect_0_sysid_0_control_slave_readdata),            //                                           .readdata
		.sysid_1_control_slave_address                    (mm_interconnect_0_sysid_1_control_slave_address),             //                      sysid_1_control_slave.address
		.sysid_1_control_slave_readdata                   (mm_interconnect_0_sysid_1_control_slave_readdata),            //                                           .readdata
		.timer_0_s1_address                               (mm_interconnect_0_timer_0_s1_address),                        //                                 timer_0_s1.address
		.timer_0_s1_write                                 (mm_interconnect_0_timer_0_s1_write),                          //                                           .write
		.timer_0_s1_readdata                              (mm_interconnect_0_timer_0_s1_readdata),                       //                                           .readdata
		.timer_0_s1_writedata                             (mm_interconnect_0_timer_0_s1_writedata),                      //                                           .writedata
		.timer_0_s1_chipselect                            (mm_interconnect_0_timer_0_s1_chipselect),                     //                                           .chipselect
		.timer_1_s1_address                               (mm_interconnect_0_timer_1_s1_address),                        //                                 timer_1_s1.address
		.timer_1_s1_write                                 (mm_interconnect_0_timer_1_s1_write),                          //                                           .write
		.timer_1_s1_readdata                              (mm_interconnect_0_timer_1_s1_readdata),                       //                                           .readdata
		.timer_1_s1_writedata                             (mm_interconnect_0_timer_1_s1_writedata),                      //                                           .writedata
		.timer_1_s1_chipselect                            (mm_interconnect_0_timer_1_s1_chipselect)                      //                                           .chipselect
	);

	MPSoC_irq_mapper irq_mapper (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.sender_irq    (cpu_0_d_irq_irq)                     //    sender.irq
	);

	MPSoC_irq_mapper_001 irq_mapper_001 (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_001_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_001_receiver1_irq),       // receiver1.irq
		.sender_irq    (cpu_1_d_irq_irq)                     //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                      // reset_in0.reset
		.reset_in1      (cpu_0_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (clk_clk),                             //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),      // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),  //          .reset_req
		.reset_req_in0  (1'b0),                                // (terminated)
		.reset_req_in1  (1'b0),                                // (terminated)
		.reset_in2      (1'b0),                                // (terminated)
		.reset_req_in2  (1'b0),                                // (terminated)
		.reset_in3      (1'b0),                                // (terminated)
		.reset_req_in3  (1'b0),                                // (terminated)
		.reset_in4      (1'b0),                                // (terminated)
		.reset_req_in4  (1'b0),                                // (terminated)
		.reset_in5      (1'b0),                                // (terminated)
		.reset_req_in5  (1'b0),                                // (terminated)
		.reset_in6      (1'b0),                                // (terminated)
		.reset_req_in6  (1'b0),                                // (terminated)
		.reset_in7      (1'b0),                                // (terminated)
		.reset_req_in7  (1'b0),                                // (terminated)
		.reset_in8      (1'b0),                                // (terminated)
		.reset_req_in8  (1'b0),                                // (terminated)
		.reset_in9      (1'b0),                                // (terminated)
		.reset_req_in9  (1'b0),                                // (terminated)
		.reset_in10     (1'b0),                                // (terminated)
		.reset_req_in10 (1'b0),                                // (terminated)
		.reset_in11     (1'b0),                                // (terminated)
		.reset_req_in11 (1'b0),                                // (terminated)
		.reset_in12     (1'b0),                                // (terminated)
		.reset_req_in12 (1'b0),                                // (terminated)
		.reset_in13     (1'b0),                                // (terminated)
		.reset_req_in13 (1'b0),                                // (terminated)
		.reset_in14     (1'b0),                                // (terminated)
		.reset_req_in14 (1'b0),                                // (terminated)
		.reset_in15     (1'b0),                                // (terminated)
		.reset_req_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (cpu_1_jtag_debug_module_reset_reset),    // reset_in1.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_002_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (cpu_1_jtag_debug_module_reset_reset),    // reset_in1.reset
		.reset_in2      (cpu_0_jtag_debug_module_reset_reset),    // reset_in2.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_003_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule

// SoC.v

// Generated using ACDS version 13.1 162 at 2025.12.20.20:41:02

`timescale 1 ps / 1 ps
module SoC (
		input  wire        clk_clk,                            //                         clk.clk
		input  wire        reset_reset_n,                      //                       reset.reset_n
		output wire [12:0] new_sdram_controller_wire_addr,     //   new_sdram_controller_wire.addr
		output wire [1:0]  new_sdram_controller_wire_ba,       //                            .ba
		output wire        new_sdram_controller_wire_cas_n,    //                            .cas_n
		output wire        new_sdram_controller_wire_cke,      //                            .cke
		output wire        new_sdram_controller_wire_cs_n,     //                            .cs_n
		inout  wire [31:0] new_sdram_controller_wire_dq,       //                            .dq
		output wire [3:0]  new_sdram_controller_wire_dqm,      //                            .dqm
		output wire        new_sdram_controller_wire_ras_n,    //                            .ras_n
		output wire        new_sdram_controller_wire_we_n,     //                            .we_n
		output wire [7:0]  led_out_external_connection_export  // led_out_external_connection.export
	);

	wire         cpu_instruction_master_waitrequest;                        // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [27:0] cpu_instruction_master_address;                            // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                               // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire  [31:0] cpu_instruction_master_readdata;                           // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire  [31:0] mm_interconnect_0_led_out_s1_writedata;                    // mm_interconnect_0:led_out_s1_writedata -> led_out:writedata
	wire   [1:0] mm_interconnect_0_led_out_s1_address;                      // mm_interconnect_0:led_out_s1_address -> led_out:address
	wire         mm_interconnect_0_led_out_s1_chipselect;                   // mm_interconnect_0:led_out_s1_chipselect -> led_out:chipselect
	wire         mm_interconnect_0_led_out_s1_write;                        // mm_interconnect_0:led_out_s1_write -> led_out:write_n
	wire  [31:0] mm_interconnect_0_led_out_s1_readdata;                     // led_out:readdata -> mm_interconnect_0:led_out_s1_readdata
	wire         cpu_data_master_waitrequest;                               // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire  [31:0] cpu_data_master_writedata;                                 // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [27:0] cpu_data_master_address;                                   // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire         cpu_data_master_write;                                     // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire         cpu_data_master_read;                                      // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire  [31:0] cpu_data_master_readdata;                                  // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_debugaccess;                               // cpu:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire   [3:0] cpu_data_master_byteenable;                                // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire   [0:0] mm_interconnect_0_sysid_control_slave_address;             // mm_interconnect_0:sysid_control_slave_address -> sysid:address
	wire  [31:0] mm_interconnect_0_sysid_control_slave_readdata;            // sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	wire         mm_interconnect_0_cpu_jtag_debug_module_waitrequest;       // cpu:jtag_debug_module_waitrequest -> mm_interconnect_0:cpu_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_cpu_jtag_debug_module_writedata;         // mm_interconnect_0:cpu_jtag_debug_module_writedata -> cpu:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_cpu_jtag_debug_module_address;           // mm_interconnect_0:cpu_jtag_debug_module_address -> cpu:jtag_debug_module_address
	wire         mm_interconnect_0_cpu_jtag_debug_module_write;             // mm_interconnect_0:cpu_jtag_debug_module_write -> cpu:jtag_debug_module_write
	wire         mm_interconnect_0_cpu_jtag_debug_module_read;              // mm_interconnect_0:cpu_jtag_debug_module_read -> cpu:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_cpu_jtag_debug_module_readdata;          // cpu:jtag_debug_module_readdata -> mm_interconnect_0:cpu_jtag_debug_module_readdata
	wire         mm_interconnect_0_cpu_jtag_debug_module_debugaccess;       // mm_interconnect_0:cpu_jtag_debug_module_debugaccess -> cpu:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_cpu_jtag_debug_module_byteenable;        // mm_interconnect_0:cpu_jtag_debug_module_byteenable -> cpu:jtag_debug_module_byteenable
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_new_sdram_controller_s1_waitrequest;     // new_sdram_controller:za_waitrequest -> mm_interconnect_0:new_sdram_controller_s1_waitrequest
	wire  [31:0] mm_interconnect_0_new_sdram_controller_s1_writedata;       // mm_interconnect_0:new_sdram_controller_s1_writedata -> new_sdram_controller:az_data
	wire  [24:0] mm_interconnect_0_new_sdram_controller_s1_address;         // mm_interconnect_0:new_sdram_controller_s1_address -> new_sdram_controller:az_addr
	wire         mm_interconnect_0_new_sdram_controller_s1_chipselect;      // mm_interconnect_0:new_sdram_controller_s1_chipselect -> new_sdram_controller:az_cs
	wire         mm_interconnect_0_new_sdram_controller_s1_write;           // mm_interconnect_0:new_sdram_controller_s1_write -> new_sdram_controller:az_wr_n
	wire         mm_interconnect_0_new_sdram_controller_s1_read;            // mm_interconnect_0:new_sdram_controller_s1_read -> new_sdram_controller:az_rd_n
	wire  [31:0] mm_interconnect_0_new_sdram_controller_s1_readdata;        // new_sdram_controller:za_data -> mm_interconnect_0:new_sdram_controller_s1_readdata
	wire         mm_interconnect_0_new_sdram_controller_s1_readdatavalid;   // new_sdram_controller:za_valid -> mm_interconnect_0:new_sdram_controller_s1_readdatavalid
	wire   [3:0] mm_interconnect_0_new_sdram_controller_s1_byteenable;      // mm_interconnect_0:new_sdram_controller_s1_byteenable -> new_sdram_controller:az_be_n
	wire  [15:0] mm_interconnect_0_timer_s1_writedata;                      // mm_interconnect_0:timer_s1_writedata -> timer:writedata
	wire   [2:0] mm_interconnect_0_timer_s1_address;                        // mm_interconnect_0:timer_s1_address -> timer:address
	wire         mm_interconnect_0_timer_s1_chipselect;                     // mm_interconnect_0:timer_s1_chipselect -> timer:chipselect
	wire         mm_interconnect_0_timer_s1_write;                          // mm_interconnect_0:timer_s1_write -> timer:write_n
	wire  [15:0] mm_interconnect_0_timer_s1_readdata;                       // timer:readdata -> mm_interconnect_0:timer_s1_readdata
	wire         irq_mapper_receiver0_irq;                                  // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                  // timer:irq -> irq_mapper:receiver1_irq
	wire  [31:0] cpu_d_irq_irq;                                             // irq_mapper:sender_irq -> cpu:d_irq
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [jtag_uart:rst_n, led_out:reset_n, mm_interconnect_0:new_sdram_controller_reset_reset_bridge_in_reset_reset, new_sdram_controller:reset_n, sysid:reset_n, timer:reset_n]
	wire         cpu_jtag_debug_module_reset_reset;                         // cpu:jtag_debug_module_resetrequest -> rst_controller:reset_in1
	wire         rst_controller_001_reset_out_reset;                        // rst_controller_001:reset_out -> [cpu:reset_n, irq_mapper:reset, mm_interconnect_0:cpu_reset_n_reset_bridge_in_reset_reset]
	wire         rst_controller_001_reset_out_reset_req;                    // rst_controller_001:reset_req -> [cpu:reset_req, rst_translator:reset_req_in]

	SoC_new_sdram_controller new_sdram_controller (
		.clk            (clk_clk),                                                 //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),                         // reset.reset_n
		.az_addr        (mm_interconnect_0_new_sdram_controller_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_new_sdram_controller_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_new_sdram_controller_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_new_sdram_controller_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_new_sdram_controller_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_new_sdram_controller_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_new_sdram_controller_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_new_sdram_controller_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_new_sdram_controller_s1_waitrequest),   //      .waitrequest
		.zs_addr        (new_sdram_controller_wire_addr),                          //  wire.export
		.zs_ba          (new_sdram_controller_wire_ba),                            //      .export
		.zs_cas_n       (new_sdram_controller_wire_cas_n),                         //      .export
		.zs_cke         (new_sdram_controller_wire_cke),                           //      .export
		.zs_cs_n        (new_sdram_controller_wire_cs_n),                          //      .export
		.zs_dq          (new_sdram_controller_wire_dq),                            //      .export
		.zs_dqm         (new_sdram_controller_wire_dqm),                           //      .export
		.zs_ras_n       (new_sdram_controller_wire_ras_n),                         //      .export
		.zs_we_n        (new_sdram_controller_wire_we_n)                           //      .export
	);

	SoC_cpu cpu (
		.clk                                   (clk_clk),                                             //                       clk.clk
		.reset_n                               (~rst_controller_001_reset_out_reset),                 //                   reset_n.reset_n
		.reset_req                             (rst_controller_001_reset_out_reset_req),              //                          .reset_req
		.d_address                             (cpu_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpu_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpu_data_master_read),                                //                          .read
		.d_readdata                            (cpu_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpu_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpu_data_master_write),                               //                          .write
		.d_writedata                           (cpu_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpu_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpu_instruction_master_read),                         //                          .read
		.i_readdata                            (cpu_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpu_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (cpu_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_cpu_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_cpu_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_cpu_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_cpu_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_cpu_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_cpu_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_cpu_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_cpu_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                     // custom_instruction_master.readra
	);

	SoC_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	SoC_timer timer (
		.clk        (clk_clk),                               //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)               //   irq.irq
	);

	SoC_sysid sysid (
		.clock    (clk_clk),                                        //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_control_slave_address)   //              .address
	);

	SoC_led_out led_out (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_led_out_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_out_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_out_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_out_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_out_s1_readdata),   //                    .readdata
		.out_port   (led_out_external_connection_export)       // external_connection.export
	);

	SoC_mm_interconnect_0 mm_interconnect_0 (
		.clock_clk_clk                                          (clk_clk),                                                   //                                        clock_clk.clk
		.cpu_reset_n_reset_bridge_in_reset_reset                (rst_controller_001_reset_out_reset),                        //                cpu_reset_n_reset_bridge_in_reset.reset
		.new_sdram_controller_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                            // new_sdram_controller_reset_reset_bridge_in_reset.reset
		.cpu_data_master_address                                (cpu_data_master_address),                                   //                                  cpu_data_master.address
		.cpu_data_master_waitrequest                            (cpu_data_master_waitrequest),                               //                                                 .waitrequest
		.cpu_data_master_byteenable                             (cpu_data_master_byteenable),                                //                                                 .byteenable
		.cpu_data_master_read                                   (cpu_data_master_read),                                      //                                                 .read
		.cpu_data_master_readdata                               (cpu_data_master_readdata),                                  //                                                 .readdata
		.cpu_data_master_write                                  (cpu_data_master_write),                                     //                                                 .write
		.cpu_data_master_writedata                              (cpu_data_master_writedata),                                 //                                                 .writedata
		.cpu_data_master_debugaccess                            (cpu_data_master_debugaccess),                               //                                                 .debugaccess
		.cpu_instruction_master_address                         (cpu_instruction_master_address),                            //                           cpu_instruction_master.address
		.cpu_instruction_master_waitrequest                     (cpu_instruction_master_waitrequest),                        //                                                 .waitrequest
		.cpu_instruction_master_read                            (cpu_instruction_master_read),                               //                                                 .read
		.cpu_instruction_master_readdata                        (cpu_instruction_master_readdata),                           //                                                 .readdata
		.cpu_jtag_debug_module_address                          (mm_interconnect_0_cpu_jtag_debug_module_address),           //                            cpu_jtag_debug_module.address
		.cpu_jtag_debug_module_write                            (mm_interconnect_0_cpu_jtag_debug_module_write),             //                                                 .write
		.cpu_jtag_debug_module_read                             (mm_interconnect_0_cpu_jtag_debug_module_read),              //                                                 .read
		.cpu_jtag_debug_module_readdata                         (mm_interconnect_0_cpu_jtag_debug_module_readdata),          //                                                 .readdata
		.cpu_jtag_debug_module_writedata                        (mm_interconnect_0_cpu_jtag_debug_module_writedata),         //                                                 .writedata
		.cpu_jtag_debug_module_byteenable                       (mm_interconnect_0_cpu_jtag_debug_module_byteenable),        //                                                 .byteenable
		.cpu_jtag_debug_module_waitrequest                      (mm_interconnect_0_cpu_jtag_debug_module_waitrequest),       //                                                 .waitrequest
		.cpu_jtag_debug_module_debugaccess                      (mm_interconnect_0_cpu_jtag_debug_module_debugaccess),       //                                                 .debugaccess
		.jtag_uart_avalon_jtag_slave_address                    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                      jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                                 .write
		.jtag_uart_avalon_jtag_slave_read                       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                                 .read
		.jtag_uart_avalon_jtag_slave_readdata                   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                                 .readdata
		.jtag_uart_avalon_jtag_slave_writedata                  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                                 .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest                (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                                 .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                 (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                                 .chipselect
		.led_out_s1_address                                     (mm_interconnect_0_led_out_s1_address),                      //                                       led_out_s1.address
		.led_out_s1_write                                       (mm_interconnect_0_led_out_s1_write),                        //                                                 .write
		.led_out_s1_readdata                                    (mm_interconnect_0_led_out_s1_readdata),                     //                                                 .readdata
		.led_out_s1_writedata                                   (mm_interconnect_0_led_out_s1_writedata),                    //                                                 .writedata
		.led_out_s1_chipselect                                  (mm_interconnect_0_led_out_s1_chipselect),                   //                                                 .chipselect
		.new_sdram_controller_s1_address                        (mm_interconnect_0_new_sdram_controller_s1_address),         //                          new_sdram_controller_s1.address
		.new_sdram_controller_s1_write                          (mm_interconnect_0_new_sdram_controller_s1_write),           //                                                 .write
		.new_sdram_controller_s1_read                           (mm_interconnect_0_new_sdram_controller_s1_read),            //                                                 .read
		.new_sdram_controller_s1_readdata                       (mm_interconnect_0_new_sdram_controller_s1_readdata),        //                                                 .readdata
		.new_sdram_controller_s1_writedata                      (mm_interconnect_0_new_sdram_controller_s1_writedata),       //                                                 .writedata
		.new_sdram_controller_s1_byteenable                     (mm_interconnect_0_new_sdram_controller_s1_byteenable),      //                                                 .byteenable
		.new_sdram_controller_s1_readdatavalid                  (mm_interconnect_0_new_sdram_controller_s1_readdatavalid),   //                                                 .readdatavalid
		.new_sdram_controller_s1_waitrequest                    (mm_interconnect_0_new_sdram_controller_s1_waitrequest),     //                                                 .waitrequest
		.new_sdram_controller_s1_chipselect                     (mm_interconnect_0_new_sdram_controller_s1_chipselect),      //                                                 .chipselect
		.sysid_control_slave_address                            (mm_interconnect_0_sysid_control_slave_address),             //                              sysid_control_slave.address
		.sysid_control_slave_readdata                           (mm_interconnect_0_sysid_control_slave_readdata),            //                                                 .readdata
		.timer_s1_address                                       (mm_interconnect_0_timer_s1_address),                        //                                         timer_s1.address
		.timer_s1_write                                         (mm_interconnect_0_timer_s1_write),                          //                                                 .write
		.timer_s1_readdata                                      (mm_interconnect_0_timer_s1_readdata),                       //                                                 .readdata
		.timer_s1_writedata                                     (mm_interconnect_0_timer_s1_writedata),                      //                                                 .writedata
		.timer_s1_chipselect                                    (mm_interconnect_0_timer_s1_chipselect)                      //                                                 .chipselect
	);

	SoC_irq_mapper irq_mapper (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.sender_irq    (cpu_d_irq_irq)                       //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                    // reset_in0.reset
		.reset_in1      (cpu_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (clk_clk),                           //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),    // reset_out.reset
		.reset_req      (),                                  // (terminated)
		.reset_req_in0  (1'b0),                              // (terminated)
		.reset_req_in1  (1'b0),                              // (terminated)
		.reset_in2      (1'b0),                              // (terminated)
		.reset_req_in2  (1'b0),                              // (terminated)
		.reset_in3      (1'b0),                              // (terminated)
		.reset_req_in3  (1'b0),                              // (terminated)
		.reset_in4      (1'b0),                              // (terminated)
		.reset_req_in4  (1'b0),                              // (terminated)
		.reset_in5      (1'b0),                              // (terminated)
		.reset_req_in5  (1'b0),                              // (terminated)
		.reset_in6      (1'b0),                              // (terminated)
		.reset_req_in6  (1'b0),                              // (terminated)
		.reset_in7      (1'b0),                              // (terminated)
		.reset_req_in7  (1'b0),                              // (terminated)
		.reset_in8      (1'b0),                              // (terminated)
		.reset_req_in8  (1'b0),                              // (terminated)
		.reset_in9      (1'b0),                              // (terminated)
		.reset_req_in9  (1'b0),                              // (terminated)
		.reset_in10     (1'b0),                              // (terminated)
		.reset_req_in10 (1'b0),                              // (terminated)
		.reset_in11     (1'b0),                              // (terminated)
		.reset_req_in11 (1'b0),                              // (terminated)
		.reset_in12     (1'b0),                              // (terminated)
		.reset_req_in12 (1'b0),                              // (terminated)
		.reset_in13     (1'b0),                              // (terminated)
		.reset_req_in13 (1'b0),                              // (terminated)
		.reset_in14     (1'b0),                              // (terminated)
		.reset_req_in14 (1'b0),                              // (terminated)
		.reset_in15     (1'b0),                              // (terminated)
		.reset_req_in15 (1'b0)                               // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
